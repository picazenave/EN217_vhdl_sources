----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08.02.2023 15:29:34
-- Design Name: 
-- Module Name: graphic_memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY graphic_memory IS
    PORT(
        clk                : IN  STD_LOGIC;
        ce                 : IN  STD_LOGIC;
        rw                 : IN  STD_LOGIC; --R/=0 W=1
        address_read_only  : IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
        address            : IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
        input              : IN  STD_LOGIC_VECTOR(47 DOWNTO 0);
        data_out_read_only : OUT STD_LOGIC_VECTOR(47 DOWNTO 0);
        data_out           : OUT STD_LOGIC_VECTOR(47 DOWNTO 0));
END graphic_memory;

ARCHITECTURE Behavioral OF graphic_memory IS
    TYPE memory_array IS ARRAY (INTEGER RANGE 0 TO 4095) OF STD_LOGIC_VECTOR(47 DOWNTO 0);
    SIGNAL memory_data : memory_array := ( --x/y
        x"100000e028f6",                --debut phrase EN217
        x"1000017028fc",
        x"100000202902",
        x"100000102908",
        x"10000070290e",
        x"100002402914",
        x"10000190291a",
        x"100001b02920",
        x"100001802926",
        x"100000c0292c",
        x"100000e02932",
        x"100001c02938",
        x"100001c0293e",
        x"100000e02944",
        x"100001e0294a",
        x"100001b02950",
        x"100002402956",
        x"10000030295c",
        x"100000202962",
        x"100000b02968",
        x"10000120296e",
        x"100001d02974",
        x"100001c0297a",
        x"100002402980",
        x"100001902986",
        x"10000180298c",
        x"100001e02992",
        x"100001b02998",
        x"10000240299e",
        x"1000015029a4",
        x"100000e029aa",
        x"1000024029b0",
        x"100000c029b6",
        x"100000a029bc",
        x"1000015029c2",
        x"100000c029c8",
        x"100001e029ce",
        x"1000015029d4",
        x"1000024029da",
        x"100000d029e0",
        x"100000e029e6",
        x"1000024029ec",
        x"1000017029f2",
        x"1000018029f8",
        x"1000016029fe",
        x"100000b02a04",
        x"100001b02a0a",
        x"100000e02a10",
        x"100001c02a16",
        x"100002402a1c",
        x"100001902a22",
        x"100001b02a28",
        x"100000e02a2e",
        x"100001602a34",
        x"100001202a3a",
        x"100000e02a40",
        x"100001b02a46",
        x"100001c02a4c",                --fin phrase EN217             
        x"0c3b89f3b89d",                --debut bongo cat
        x"0c3bca03bc9c",
        x"0c3c0a13c09c",
        x"0c3c4a23c49b",
        x"0c3c8a33c89a",
        x"0c3cca43cc99",
        x"0c3d0a53d099",
        x"0c3d4a63d498",
        x"0c3d8a73d897",
        x"0c3dca83dc96",
        x"0c3e0a93e095",
        x"0c3e4aa3e495",
        x"0c3e8ab3e894",
        x"0c3ecab3ec93",
        x"0c3f0ac3f092",
        x"0c3f4ad3f492",
        x"0c3f8ae3f892",
        x"0c3fcb13fc91",
        x"0c400b340090",
        x"0c404b64048f",
        x"0c408b94088e",
        x"0c40cbc40c8a",
        x"0c410bf41086",
        x"0c414c141483",
        x"0c418c341880",
        x"0c41cc541c7d",
        x"0c420c74207b",
        x"0c424c842479",
        x"0c428ca42876",
        x"0c42ccc42c74",
        x"0c430ce43071",
        x"0c434cf4346f",
        x"0c438d14386c",
        x"0c43cd243c69",
        x"0c440d444066",
        x"0c444d544463",
        x"0c448d644860",
        x"0c44cd844c5e",
        x"0c450d94505b",
        x"0c454db45459",
        x"0c458dc45857",
        x"0c45cdd45c54",
        x"0c460df46053",
        x"0c464e046451",
        x"0c468e14684f",
        x"0c46ce246c4d",
        x"0c470e34704c",
        x"0c4741f4741e",
        x"0c474e54744a",
        x"0c478214781e",
        x"0c478e647848",
        x"0c47c2447c1e",
        x"0c47ce747c46",
        x"0c480264801e",
        x"0c480e848045",
        x"0c484294841e",
        x"0c484e948443",
        x"0c4882b4881e",
        x"0c488ea48841",
        x"0c48c2e48c1e",
        x"0c48ceb48c3f",
        x"0c490304901e",
        x"0c490ec4903c",
        x"0c494324941e",
        x"0c494ee4943a",
        x"0c498354981e",
        x"0c498ef49838",
        x"0c49cf049c1e",
        x"0c4a0f14a01e",
        x"0c4a4f24a41e",
        x"0c4a8f44a81e",
        x"0c4acf44ac1e",
        x"0c4b0f54b01e",
        x"0c4b4bd4b41e",
        x"0c4b4f64b4c4",
        x"0c4b8bc4b81e",
        x"0c4b8f74b8c5",
        x"0c4bcbb4bc1e",
        x"0c4bcf94bcc6",
        x"0c4c0bb4c01f",
        x"0c4c0fa4c0c7",
        x"0c4c4ba4c41f",
        x"0c4c4fb4c4c7",
        x"0c4c8ba4c81f",
        x"0c4c8fc4c8c7",
        x"0c4ccba4cc1f",
        x"0c4ccfd4ccc7",
        x"0c4d0ba4d020",
        x"0c4d0fe4d0c7",
        x"0c4d4ba4d420",
        x"0c4d4ff4d4c7",
        x"0c4d8bb4d821",
        x"0c4d9004d8c7",
        x"0c4dcae4dc21",
        x"0c4dcbb4dcb2",
        x"0c4dd014dcc7",
        x"0c4e0ad4e021",
        x"0c4e0bc4e0b3",
        x"0c4e1024e0c7",
        x"0c4e4a04e422",
        x"0c4e4ad4e4a3",
        x"0c4e4bd4e4b3",
        x"0c4e5034e4c6",
        x"0c4e89f4e822",
        x"0c4e8ad4e8a4",
        x"0c4e8bf4e8b3",
        x"0c4e9034e8c3",
        x"0c4ec9e4ec23",
        x"0c4ecac4eca7",
        x"0c4ed044ecb3",
        x"0c4f09e4f023",
        x"0c4f1054f0b3",
        x"0c4f49e4f423",
        x"0c4f5064f4b2",
        x"0c4f89e4f823",
        x"0c4f9064f8b1",
        x"0c4fc9d4fc24",
        x"0c4fd074fcb0",
        x"0c5009c50024",
        x"0c50108500af",
        x"0c5049250424",
        x"0c50509504a3",
        x"0c5089250824",
        x"0c5090a508a2",
        x"0c50c9150c24",
        x"0c50d0a50ca1",
        x"0c5109151024",
        x"0c5110b510a0",
        x"0c5149251425",
        x"0c5150c5149f",
        x"0c5186e51825",
        x"0c5189451870",
        x"0c5190c5189c",
        x"0c51c6c51c25",
        x"0c51d0d51c73",
        x"0c5206c52025",
        x"0c5210d52074",
        x"0c5246b52426",
        x"0c5250d52475",
        x"0c5286b52826",
        x"0c5290e52876",
        x"0c52c6b52c26",
        x"0c52d0f52c77",
        x"0c5306b53027",
        x"0c5310f53077",
        x"0c5346b53427",
        x"0c5351053477",
        x"0c5386b53827",
        x"0c5391053877",
        x"0c53c6b53c26",
        x"0c53d1053c77",
        x"0c5406b54026",
        x"0c5411054077",
        x"0c5446c54425",
        x"0c544d454476",
        x"0c54510544d9",
        x"0c5486d54824",
        x"0c548d154875",
        x"0c54910548dc",
        x"0c54ccd54c23",
        x"0c54d1054cdf",
        x"0c550c855023",
        x"0c55110550e3",
        x"0c554c355422",
        x"0c55510554e7",
        x"0c558be55821",
        x"0c5590f558ea",
        x"0c55cb955c20",
        x"0c55d0e55ced",
        x"0c560b556020",
        x"0c5610d560f1",
        x"0c564b05641f",
        x"0c5650b564f3",
        x"0c568ad5681f",
        x"0c56909568f6",
        x"0c56ca956c1e",
        x"0c570a45701e",
        x"0c574a05741d",
        x"0c5789c5781d",
        x"0c57c9857c1c",
        x"0c580935801c",
        x"0c5846a5841b",
        x"0c5848f5846d",
        x"0c588695881b",
        x"0c5888b5886e",
        x"0c58c6958c1a",
        x"0c58c8758c6f",
        x"0c590695901a",
        x"0c5908359070",
        x"0c5946a5941a",
        x"0c5947e59471",
        x"0c5986b59819",
        x"0c5987a59872",
        x"0c59c6c59c19",
        x"0c59c7659c73",
        x"0c5a06d5a018",
        x"0c5a46e5a418",
        x"0c5a86e5a818",
        x"0c5ac6f5ac17",
        x"0c5b0705b017",
        x"0c5b4705b416",
        x"0c5b8715b816",
        x"0c5bc725bc16",
        x"0c5c0725c015",
        x"0c5c4735c415",
        x"0c5c8735c815",
        x"0c5cc735cc14",
        x"0c5d0735d014",
        x"0c5d42f5d413",
        x"0c5d4735d43b",
        x"0c5d82e5d813",
        x"0c5d8735d83f",
        x"0c5dc2e5dc13",
        x"0c5dc735dc43",
        x"0c5e02d5e013",
        x"0c5e0735e046",
        x"0c5e42a5e412",
        x"0c5e4735e449",
        x"0c5e8265e812",
        x"0c5e8725e84b",
        x"0c5ec235ec12",
        x"0c5ec715ec4e",
        x"0c5f01d5f012",
        x"0c5f06f5f053",
        x"0c5f4185f412",
        x"0c5f46e5f456",
        x"0c5f8145f812",
        x"0c5f86b5f859",                --fin bongo cat
        x"0c02cd302c0b",                --debut qr
        x"0c030d30300b",
        x"0c034d30340b",
        x"0c038d30380b",
        x"0c03cd303c0b",
        x"0c040d30400b",
        x"0c044d30440b",
        x"0c048d30480b",
        x"0c04c1304c0b",
        x"0c04c5e04c3f",
        x"0c04c6a04c64",
        x"0c04c7604c70",
        x"0c04c9c04c7d",
        x"0c04cd304cc7",
        x"0c050130500b",
        x"0c0505e0503f",
        x"0c0506a05064",
        x"0c0507605070",
        x"0c0509c0507d",
        x"0c050d3050c7",
        x"0c054130540b",
        x"0c0545e0543f",
        x"0c0546a05464",
        x"0c0547605470",
        x"0c0549c0547d",
        x"0c054d3054c7",
        x"0c058130580b",
        x"0c0585e0583f",
        x"0c0586a05864",
        x"0c0587605870",
        x"0c0589c0587d",
        x"0c058d3058c7",
        x"0c05c1305c0b",
        x"0c05c5e05c3f",
        x"0c05c6a05c64",
        x"0c05c7605c70",
        x"0c05c9c05c7d",
        x"0c05cd305cc7",
        x"0c060130600b",
        x"0c0605e0603f",
        x"0c0606a06064",
        x"0c0607606070",
        x"0c0609c0607d",
        x"0c060d3060c7",
        x"0c064130640b",
        x"0c0643806419",
        x"0c0644b0643f",
        x"0c0645706451",
        x"0c0647606470",
        x"0c064830647d",
        x"0c0648f06489",
        x"0c0649c06495",
        x"0c064c0064a2",
        x"0c064d3064c7",
        x"0c068130680b",
        x"0c0683806819",
        x"0c0684b0683f",
        x"0c0685706851",
        x"0c0687606870",
        x"0c068830687d",
        x"0c0688f06889",
        x"0c0689c06895",
        x"0c068c0068a2",
        x"0c068d3068c7",
        x"0c06c1306c0b",
        x"0c06c3806c19",
        x"0c06c4b06c3f",
        x"0c06c5706c51",
        x"0c06c7606c70",
        x"0c06c8306c7d",
        x"0c06c8f06c89",
        x"0c06c9c06c95",
        x"0c06cc006ca2",
        x"0c06cd306cc7",
        x"0c070130700b",
        x"0c0703807019",
        x"0c0704b0703f",
        x"0c0705707051",
        x"0c0707607070",
        x"0c070830707d",
        x"0c0708f07089",
        x"0c0709c07095",
        x"0c070c0070a2",
        x"0c070d3070c7",
        x"0c074130740b",
        x"0c0743807419",
        x"0c0744b0743f",
        x"0c0745707451",
        x"0c0747607470",
        x"0c074830747d",
        x"0c0748f07489",
        x"0c0749c07495",
        x"0c074c0074a2",
        x"0c074d3074c7",
        x"0c078130780b",
        x"0c0783807819",
        x"0c0784b0783f",
        x"0c0785707851",
        x"0c0787607870",
        x"0c078830787d",
        x"0c0788f07889",
        x"0c0789c07895",
        x"0c078c0078a2",
        x"0c078d3078c7",
        x"0c07c1307c0b",
        x"0c07c1f07c19",
        x"0c07c3807c32",
        x"0c07c4507c3f",
        x"0c07c6a07c57",
        x"0c07c9c07c7d",
        x"0c07ca807ca2",
        x"0c07cc007cbb",
        x"0c07cd307cc7",
        x"0c080130800b",
        x"0c0801f08019",
        x"0c0803808032",
        x"0c080450803f",
        x"0c0806a08057",
        x"0c0809c0807d",
        x"0c080a8080a2",
        x"0c080c0080bb",
        x"0c080d3080c7",
        x"0c084130840b",
        x"0c0841f08419",
        x"0c0843808432",
        x"0c084450843f",
        x"0c0846a08457",
        x"0c0849c0847d",
        x"0c084a8084a2",
        x"0c084c0084bb",
        x"0c084d3084c7",
        x"0c088130880b",
        x"0c0881f08819",
        x"0c0883808832",
        x"0c088450883f",
        x"0c0886a08857",
        x"0c0889c0887d",
        x"0c088a8088a2",
        x"0c088c0088bb",
        x"0c088d3088c7",
        x"0c08c1308c0b",
        x"0c08c1f08c19",
        x"0c08c3808c32",
        x"0c08c4508c3f",
        x"0c08c6a08c57",
        x"0c08c9c08c7d",
        x"0c08ca808ca2",
        x"0c08cc008cbb",
        x"0c08cd308cc7",
        x"0c090130900b",
        x"0c0901f09019",
        x"0c0903809032",
        x"0c090450903f",
        x"0c0906a09057",
        x"0c0909c0907d",
        x"0c090a8090a2",
        x"0c090c0090bb",
        x"0c090d3090c7",
        x"0c094130940b",
        x"0c0941f09419",
        x"0c0943809432",
        x"0c094510943f",
        x"0c0948309476",
        x"0c0949c09495",
        x"0c094a8094a2",
        x"0c094c0094bb",
        x"0c094d3094c7",
        x"0c098130980b",
        x"0c0981f09819",
        x"0c0983809832",
        x"0c098510983f",
        x"0c0988309876",
        x"0c0989c09895",
        x"0c098a8098a2",
        x"0c098c0098bb",
        x"0c098d3098c7",
        x"0c09c1309c0b",
        x"0c09c1f09c19",
        x"0c09c3809c32",
        x"0c09c5109c3f",
        x"0c09c8309c76",
        x"0c09c9c09c95",
        x"0c09ca809ca2",
        x"0c09cc009cbb",
        x"0c09cd309cc7",
        x"0c0a0130a00b",
        x"0c0a01f0a019",
        x"0c0a0380a032",
        x"0c0a0510a03f",
        x"0c0a0830a076",
        x"0c0a09c0a095",
        x"0c0a0a80a0a2",
        x"0c0a0c00a0bb",
        x"0c0a0d30a0c7",
        x"0c0a4130a40b",
        x"0c0a41f0a419",
        x"0c0a4380a432",
        x"0c0a4510a43f",
        x"0c0a4830a476",
        x"0c0a49c0a495",
        x"0c0a4a80a4a2",
        x"0c0a4c00a4bb",
        x"0c0a4d30a4c7",
        x"0c0a8130a80b",
        x"0c0a81f0a819",
        x"0c0a8380a832",
        x"0c0a8510a83f",
        x"0c0a8830a876",
        x"0c0a89c0a895",
        x"0c0a8a80a8a2",
        x"0c0a8c00a8bb",
        x"0c0a8d30a8c7",
        x"0c0ac130ac0b",
        x"0c0ac1f0ac19",
        x"0c0ac380ac32",
        x"0c0ac510ac3f",
        x"0c0ac830ac76",
        x"0c0ac9c0ac95",
        x"0c0aca80aca2",
        x"0c0acc00acbb",
        x"0c0acd30acc7",
        x"0c0b0130b00b",
        x"0c0b01f0b019",
        x"0c0b0380b032",
        x"0c0b0640b03f",
        x"0c0b0760b070",
        x"0c0b0890b083",
        x"0c0b09c0b08f",
        x"0c0b0a80b0a2",
        x"0c0b0c00b0bb",
        x"0c0b0d30b0c7",
        x"0c0b4130b40b",
        x"0c0b41f0b419",
        x"0c0b4380b432",
        x"0c0b4640b43f",
        x"0c0b4760b470",
        x"0c0b4890b483",
        x"0c0b49c0b48f",
        x"0c0b4a80b4a2",
        x"0c0b4c00b4bb",
        x"0c0b4d30b4c7",
        x"0c0b8130b80b",
        x"0c0b81f0b819",
        x"0c0b8380b832",
        x"0c0b8640b83f",
        x"0c0b8760b870",
        x"0c0b8890b883",
        x"0c0b89c0b88f",
        x"0c0b8a80b8a2",
        x"0c0b8c00b8bb",
        x"0c0b8d30b8c7",
        x"0c0bc130bc0b",
        x"0c0bc1f0bc19",
        x"0c0bc380bc32",
        x"0c0bc640bc3f",
        x"0c0bc760bc70",
        x"0c0bc890bc83",
        x"0c0bc9c0bc8f",
        x"0c0bca80bca2",
        x"0c0bcc00bcbb",
        x"0c0bcd30bcc7",
        x"0c0c0130c00b",
        x"0c0c01f0c019",
        x"0c0c0380c032",
        x"0c0c0640c03f",
        x"0c0c0760c070",
        x"0c0c0890c083",
        x"0c0c09c0c08f",
        x"0c0c0a80c0a2",
        x"0c0c0c00c0bb",
        x"0c0c0d30c0c7",
        x"0c0c4130c40b",
        x"0c0c41f0c419",
        x"0c0c4380c432",
        x"0c0c4640c43f",
        x"0c0c4760c470",
        x"0c0c4890c483",
        x"0c0c49c0c48f",
        x"0c0c4a80c4a2",
        x"0c0c4c00c4bb",
        x"0c0c4d30c4c7",
        x"0c0c8130c80b",
        x"0c0c8380c819",
        x"0c0c8450c83f",
        x"0c0c8570c84b",
        x"0c0c8890c876",
        x"0c0c89c0c895",
        x"0c0c8c00c8a2",
        x"0c0c8d30c8c7",
        x"0c0cc130cc0b",
        x"0c0cc380cc19",
        x"0c0cc450cc3f",
        x"0c0cc570cc4b",
        x"0c0cc890cc76",
        x"0c0cc9c0cc95",
        x"0c0ccc00cca2",
        x"0c0ccd30ccc7",
        x"0c0d0130d00b",
        x"0c0d0380d019",
        x"0c0d0450d03f",
        x"0c0d0570d04b",
        x"0c0d0890d076",
        x"0c0d09c0d095",
        x"0c0d0c00d0a2",
        x"0c0d0d30d0c7",
        x"0c0d4130d40b",
        x"0c0d4380d419",
        x"0c0d4450d43f",
        x"0c0d4570d44b",
        x"0c0d4890d476",
        x"0c0d49c0d495",
        x"0c0d4c00d4a2",
        x"0c0d4d30d4c7",
        x"0c0d8130d80b",
        x"0c0d8380d819",
        x"0c0d8450d83f",
        x"0c0d8570d84b",
        x"0c0d8890d876",
        x"0c0d89c0d895",
        x"0c0d8c00d8a2",
        x"0c0d8d30d8c7",
        x"0c0dc130dc0b",
        x"0c0dc380dc19",
        x"0c0dc450dc3f",
        x"0c0dc570dc4b",
        x"0c0dc890dc76",
        x"0c0dc9c0dc95",
        x"0c0dcc00dca2",
        x"0c0dcd30dcc7",
        x"0c0e0130e00b",
        x"0c0e0450e03f",
        x"0c0e0510e04b",
        x"0c0e05e0e057",
        x"0c0e06a0e064",
        x"0c0e0760e070",
        x"0c0e0830e07d",
        x"0c0e08f0e089",
        x"0c0e09c0e095",
        x"0c0e0d30e0c7",
        x"0c0e4130e40b",
        x"0c0e4450e43f",
        x"0c0e4510e44b",
        x"0c0e45e0e457",
        x"0c0e46a0e464",
        x"0c0e4760e470",
        x"0c0e4830e47d",
        x"0c0e48f0e489",
        x"0c0e49c0e495",
        x"0c0e4d30e4c7",
        x"0c0e8130e80b",
        x"0c0e8450e83f",
        x"0c0e8510e84b",
        x"0c0e85e0e857",
        x"0c0e86a0e864",
        x"0c0e8760e870",
        x"0c0e8830e87d",
        x"0c0e88f0e889",
        x"0c0e89c0e895",
        x"0c0e8d30e8c7",
        x"0c0ec130ec0b",
        x"0c0ec450ec3f",
        x"0c0ec510ec4b",
        x"0c0ec5e0ec57",
        x"0c0ec6a0ec64",
        x"0c0ec760ec70",
        x"0c0ec830ec7d",
        x"0c0ec8f0ec89",
        x"0c0ec9c0ec95",
        x"0c0ecd30ecc7",
        x"0c0f0130f00b",
        x"0c0f0450f03f",
        x"0c0f0510f04b",
        x"0c0f05e0f057",
        x"0c0f06a0f064",
        x"0c0f0760f070",
        x"0c0f0830f07d",
        x"0c0f08f0f089",
        x"0c0f09c0f095",
        x"0c0f0d30f0c7",
        x"0c0f4130f40b",
        x"0c0f4450f43f",
        x"0c0f4510f44b",
        x"0c0f45e0f457",
        x"0c0f46a0f464",
        x"0c0f4760f470",
        x"0c0f4830f47d",
        x"0c0f48f0f489",
        x"0c0f49c0f495",
        x"0c0f4d30f4c7",
        x"0c0f8450f80b",
        x"0c0f86a0f857",
        x"0c0f87d0f870",
        x"0c0f8d30f88f",
        x"0c0fc450fc0b",
        x"0c0fc6a0fc57",
        x"0c0fc7d0fc70",
        x"0c0fcd30fc8f",
        x"0c100451000b",
        x"0c1006a10057",
        x"0c1007d10070",
        x"0c100d31008f",
        x"0c104451040b",
        x"0c1046a10457",
        x"0c1047d10470",
        x"0c104d31048f",
        x"0c108451080b",
        x"0c1086a10857",
        x"0c1087d10870",
        x"0c108d31088f",
        x"0c10c4510c0b",
        x"0c10c6a10c57",
        x"0c10c7d10c70",
        x"0c10cd310c8f",
        x"0c110191100b",
        x"0c110261101f",
        x"0c110321102c",
        x"0c1103e11038",
        x"0c110511104b",
        x"0c1106411057",
        x"0c1108911076",
        x"0c110a8110a2",
        x"0c110d3110c7",
        x"0c114191140b",
        x"0c114261141f",
        x"0c114321142c",
        x"0c1143e11438",
        x"0c114511144b",
        x"0c1146411457",
        x"0c1148911476",
        x"0c114a8114a2",
        x"0c114d3114c7",
        x"0c118191180b",
        x"0c118261181f",
        x"0c118321182c",
        x"0c1183e11838",
        x"0c118511184b",
        x"0c1186411857",
        x"0c1188911876",
        x"0c118a8118a2",
        x"0c118d3118c7",
        x"0c11c1911c0b",
        x"0c11c2611c1f",
        x"0c11c3211c2c",
        x"0c11c3e11c38",
        x"0c11c5111c4b",
        x"0c11c6411c57",
        x"0c11c8911c76",
        x"0c11ca811ca2",
        x"0c11cd311cc7",
        x"0c120191200b",
        x"0c120261201f",
        x"0c120321202c",
        x"0c1203e12038",
        x"0c120511204b",
        x"0c1206412057",
        x"0c1208912076",
        x"0c120a8120a2",
        x"0c120d3120c7",
        x"0c124191240b",
        x"0c124261241f",
        x"0c124321242c",
        x"0c1243e12438",
        x"0c124511244b",
        x"0c1246412457",
        x"0c1248912476",
        x"0c124a8124a2",
        x"0c124d3124c7",
        x"0c128191280b",
        x"0c128261281f",
        x"0c1283e12838",
        x"0c1288312851",
        x"0c1289512889",
        x"0c128a21289c",
        x"0c128ae128a8",
        x"0c128bb128b5",
        x"0c128d3128c7",
        x"0c12c1912c0b",
        x"0c12c2612c1f",
        x"0c12c3e12c38",
        x"0c12c8312c51",
        x"0c12c9512c89",
        x"0c12ca212c9c",
        x"0c12cae12ca8",
        x"0c12cbb12cb5",
        x"0c12cd312cc7",
        x"0c130191300b",
        x"0c130261301f",
        x"0c1303e13038",
        x"0c1308313051",
        x"0c1309513089",
        x"0c130a21309c",
        x"0c130ae130a8",
        x"0c130bb130b5",
        x"0c130d3130c7",
        x"0c134191340b",
        x"0c134261341f",
        x"0c1343e13438",
        x"0c1348313451",
        x"0c1349513489",
        x"0c134a21349c",
        x"0c134ae134a8",
        x"0c134bb134b5",
        x"0c134d3134c7",
        x"0c138191380b",
        x"0c138261381f",
        x"0c1383e13838",
        x"0c1388313851",
        x"0c1389513889",
        x"0c138a21389c",
        x"0c138ae138a8",
        x"0c138bb138b5",
        x"0c138d3138c7",
        x"0c13c1913c0b",
        x"0c13c2613c1f",
        x"0c13c3e13c38",
        x"0c13c8313c51",
        x"0c13c9513c89",
        x"0c13ca213c9c",
        x"0c13cae13ca8",
        x"0c13cbb13cb5",
        x"0c13cd313cc7",
        x"0c140191400b",
        x"0c140261401f",
        x"0c1403e14038",
        x"0c1408314051",
        x"0c1409514089",
        x"0c140a21409c",
        x"0c140ae140a8",
        x"0c140bb140b5",
        x"0c140d3140c7",
        x"0c1441f1440b",
        x"0c144321442c",
        x"0c1444b14438",
        x"0c1445714451",
        x"0c144831447d",
        x"0c1449514489",
        x"0c144a8144a2",
        x"0c144bb144ae",
        x"0c144d3144c1",
        x"0c1481f1480b",
        x"0c148321482c",
        x"0c1484b14838",
        x"0c1485714851",
        x"0c148831487d",
        x"0c1489514889",
        x"0c148a8148a2",
        x"0c148bb148ae",
        x"0c148d3148c1",
        x"0c14c1f14c0b",
        x"0c14c3214c2c",
        x"0c14c4b14c38",
        x"0c14c5714c51",
        x"0c14c8314c7d",
        x"0c14c9514c89",
        x"0c14ca814ca2",
        x"0c14cbb14cae",
        x"0c14cd314cc1",
        x"0c1501f1500b",
        x"0c150321502c",
        x"0c1504b15038",
        x"0c1505715051",
        x"0c150831507d",
        x"0c1509515089",
        x"0c150a8150a2",
        x"0c150bb150ae",
        x"0c150d3150c1",
        x"0c1541f1540b",
        x"0c154321542c",
        x"0c1544b15438",
        x"0c1545715451",
        x"0c154831547d",
        x"0c1549515489",
        x"0c154a8154a2",
        x"0c154bb154ae",
        x"0c154d3154c1",
        x"0c1581f1580b",
        x"0c158321582c",
        x"0c1584b15838",
        x"0c1585715851",
        x"0c158831587d",
        x"0c1589515889",
        x"0c158a8158a2",
        x"0c158bb158ae",
        x"0c158d3158c1",
        x"0c15c1315c0b",
        x"0c15c2615c19",
        x"0c15c4b15c45",
        x"0c15c5715c51",
        x"0c15c7015c5e",
        x"0c15c7d15c76",
        x"0c15c9515c83",
        x"0c15ca815c9c",
        x"0c15cc115cbb",
        x"0c15cd315cc7",
        x"0c160131600b",
        x"0c1602616019",
        x"0c1604b16045",
        x"0c1605716051",
        x"0c160701605e",
        x"0c1607d16076",
        x"0c1609516083",
        x"0c160a81609c",
        x"0c160c1160bb",
        x"0c160d3160c7",
        x"0c164131640b",
        x"0c1642616419",
        x"0c1644b16445",
        x"0c1645716451",
        x"0c164701645e",
        x"0c1647d16476",
        x"0c1649516483",
        x"0c164a81649c",
        x"0c164c1164bb",
        x"0c164d3164c7",
        x"0c168131680b",
        x"0c1682616819",
        x"0c1684b16845",
        x"0c1685716851",
        x"0c168701685e",
        x"0c1687d16876",
        x"0c1689516883",
        x"0c168a81689c",
        x"0c168c1168bb",
        x"0c168d3168c7",
        x"0c16c1316c0b",
        x"0c16c2616c19",
        x"0c16c4b16c45",
        x"0c16c5716c51",
        x"0c16c7016c5e",
        x"0c16c7d16c76",
        x"0c16c9516c83",
        x"0c16ca816c9c",
        x"0c16cc116cbb",
        x"0c16cd316cc7",
        x"0c170131700b",
        x"0c1702617019",
        x"0c1704b17045",
        x"0c1705717051",
        x"0c170701705e",
        x"0c1707d17076",
        x"0c1709517083",
        x"0c170a81709c",
        x"0c170c1170bb",
        x"0c170d3170c7",
        x"0c1742c1740b",
        x"0c174511744b",
        x"0c174641745e",
        x"0c174831746a",
        x"0c174b5174a2",
        x"0c174d3174c1",
        x"0c1782c1780b",
        x"0c178511784b",
        x"0c178641785e",
        x"0c178831786a",
        x"0c178b5178a2",
        x"0c178d3178c1",
        x"0c17c2c17c0b",
        x"0c17c5117c4b",
        x"0c17c6417c5e",
        x"0c17c8317c6a",
        x"0c17cb517ca2",
        x"0c17cd317cc1",
        x"0c1802c1800b",
        x"0c180511804b",
        x"0c180641805e",
        x"0c180831806a",
        x"0c180b5180a2",
        x"0c180d3180c1",
        x"0c1842c1840b",
        x"0c184511844b",
        x"0c184641845e",
        x"0c184831846a",
        x"0c184b5184a2",
        x"0c184d3184c1",
        x"0c1882c1880b",
        x"0c188511884b",
        x"0c188641885e",
        x"0c188831886a",
        x"0c188b5188a2",
        x"0c188d3188c1",
        x"0c18c1918c0b",
        x"0c18c2618c1f",
        x"0c18c3e18c2c",
        x"0c18c5118c4b",
        x"0c18c5e18c57",
        x"0c18c7618c64",
        x"0c18c8f18c83",
        x"0c18ca218c95",
        x"0c18cbb18cae",
        x"0c18cd318cc7",
        x"0c190191900b",
        x"0c190261901f",
        x"0c1903e1902c",
        x"0c190511904b",
        x"0c1905e19057",
        x"0c1907619064",
        x"0c1908f19083",
        x"0c190a219095",
        x"0c190bb190ae",
        x"0c190d3190c7",
        x"0c194191940b",
        x"0c194261941f",
        x"0c1943e1942c",
        x"0c194511944b",
        x"0c1945e19457",
        x"0c1947619464",
        x"0c1948f19483",
        x"0c194a219495",
        x"0c194bb194ae",
        x"0c194d3194c7",
        x"0c198191980b",
        x"0c198261981f",
        x"0c1983e1982c",
        x"0c198511984b",
        x"0c1985e19857",
        x"0c1987619864",
        x"0c1988f19883",
        x"0c198a219895",
        x"0c198bb198ae",
        x"0c198d3198c7",
        x"0c19c1919c0b",
        x"0c19c2619c1f",
        x"0c19c3e19c2c",
        x"0c19c5119c4b",
        x"0c19c5e19c57",
        x"0c19c7619c64",
        x"0c19c8f19c83",
        x"0c19ca219c95",
        x"0c19cbb19cae",
        x"0c19cd319cc7",
        x"0c1a0191a00b",
        x"0c1a0261a01f",
        x"0c1a03e1a02c",
        x"0c1a0511a04b",
        x"0c1a05e1a057",
        x"0c1a0761a064",
        x"0c1a08f1a083",
        x"0c1a0a21a095",
        x"0c1a0bb1a0ae",
        x"0c1a0d31a0c7",
        x"0c1a4131a40b",
        x"0c1a44b1a42c",
        x"0c1a4571a451",
        x"0c1a46a1a45e",
        x"0c1a4831a47d",
        x"0c1a49c1a495",
        x"0c1a4d31a4c7",
        x"0c1a8131a80b",
        x"0c1a84b1a82c",
        x"0c1a8571a851",
        x"0c1a86a1a85e",
        x"0c1a8831a87d",
        x"0c1a89c1a895",
        x"0c1a8d31a8c7",
        x"0c1ac131ac0b",
        x"0c1ac4b1ac2c",
        x"0c1ac571ac51",
        x"0c1ac6a1ac5e",
        x"0c1ac831ac7d",
        x"0c1ac9c1ac95",
        x"0c1acd31acc7",
        x"0c1b0131b00b",
        x"0c1b04b1b02c",
        x"0c1b0571b051",
        x"0c1b06a1b05e",
        x"0c1b0831b07d",
        x"0c1b09c1b095",
        x"0c1b0d31b0c7",
        x"0c1b4131b40b",
        x"0c1b44b1b42c",
        x"0c1b4571b451",
        x"0c1b46a1b45e",
        x"0c1b4831b47d",
        x"0c1b49c1b495",
        x"0c1b4d31b4c7",
        x"0c1b8131b80b",
        x"0c1b84b1b82c",
        x"0c1b8571b851",
        x"0c1b86a1b85e",
        x"0c1b8831b87d",
        x"0c1b89c1b895",
        x"0c1b8d31b8c7",
        x"0c1bc131bc0b",
        x"0c1bc4b1bc2c",
        x"0c1bc571bc51",
        x"0c1bc6a1bc5e",
        x"0c1bc831bc7d",
        x"0c1bc9c1bc95",
        x"0c1bcd31bcc7",
        x"0c1c0131c00b",
        x"0c1c02c1c01f",
        x"0c1c0451c03e",
        x"0c1c05e1c057",
        x"0c1c07d1c06a",
        x"0c1c0891c083",
        x"0c1c0a21c09c",
        x"0c1c0bb1c0a8",
        x"0c1c0d31c0c1",
        x"0c1c4131c40b",
        x"0c1c42c1c41f",
        x"0c1c4451c43e",
        x"0c1c45e1c457",
        x"0c1c47d1c46a",
        x"0c1c4891c483",
        x"0c1c4a21c49c",
        x"0c1c4bb1c4a8",
        x"0c1c4d31c4c1",
        x"0c1c8131c80b",
        x"0c1c82c1c81f",
        x"0c1c8451c83e",
        x"0c1c85e1c857",
        x"0c1c87d1c86a",
        x"0c1c8891c883",
        x"0c1c8a21c89c",
        x"0c1c8bb1c8a8",
        x"0c1c8d31c8c1",
        x"0c1cc131cc0b",
        x"0c1cc2c1cc1f",
        x"0c1cc451cc3e",
        x"0c1cc5e1cc57",
        x"0c1cc7d1cc6a",
        x"0c1cc891cc83",
        x"0c1cca21cc9c",
        x"0c1ccbb1cca8",
        x"0c1ccd31ccc1",
        x"0c1d0131d00b",
        x"0c1d02c1d01f",
        x"0c1d0451d03e",
        x"0c1d05e1d057",
        x"0c1d07d1d06a",
        x"0c1d0891d083",
        x"0c1d0a21d09c",
        x"0c1d0bb1d0a8",
        x"0c1d0d31d0c1",
        x"0c1d4131d40b",
        x"0c1d42c1d41f",
        x"0c1d4451d43e",
        x"0c1d45e1d457",
        x"0c1d47d1d46a",
        x"0c1d4891d483",
        x"0c1d4a21d49c",
        x"0c1d4bb1d4a8",
        x"0c1d4d31d4c1",
        x"0c1d8321d80b",
        x"0c1d8451d838",
        x"0c1d85e1d84b",
        x"0c1d8761d870",
        x"0c1d8831d87d",
        x"0c1d8951d889",
        x"0c1d8d31d8ae",
        x"0c1dc321dc0b",
        x"0c1dc451dc38",
        x"0c1dc5e1dc4b",
        x"0c1dc761dc70",
        x"0c1dc831dc7d",
        x"0c1dc951dc89",
        x"0c1dcd31dcae",
        x"0c1e0321e00b",
        x"0c1e0451e038",
        x"0c1e05e1e04b",
        x"0c1e0761e070",
        x"0c1e0831e07d",
        x"0c1e0951e089",
        x"0c1e0d31e0ae",
        x"0c1e4321e40b",
        x"0c1e4451e438",
        x"0c1e45e1e44b",
        x"0c1e4761e470",
        x"0c1e4831e47d",
        x"0c1e4951e489",
        x"0c1e4d31e4ae",
        x"0c1e8321e80b",
        x"0c1e8451e838",
        x"0c1e85e1e84b",
        x"0c1e8761e870",
        x"0c1e8831e87d",
        x"0c1e8951e889",
        x"0c1e8d31e8ae",
        x"0c1ec321ec0b",
        x"0c1ec451ec38",
        x"0c1ec5e1ec4b",
        x"0c1ec761ec70",
        x"0c1ec831ec7d",
        x"0c1ec951ec89",
        x"0c1ecd31ecae",
        x"0c1f0191f00b",
        x"0c1f0261f01f",
        x"0c1f0451f038",
        x"0c1f05e1f051",
        x"0c1f0761f06a",
        x"0c1f0b51f083",
        x"0c1f0d31f0c7",
        x"0c1f4191f40b",
        x"0c1f4261f41f",
        x"0c1f4451f438",
        x"0c1f45e1f451",
        x"0c1f4761f46a",
        x"0c1f4b51f483",
        x"0c1f4d31f4c7",
        x"0c1f8191f80b",
        x"0c1f8261f81f",
        x"0c1f8451f838",
        x"0c1f85e1f851",
        x"0c1f8761f86a",
        x"0c1f8b51f883",
        x"0c1f8d31f8c7",
        x"0c1fc191fc0b",
        x"0c1fc261fc1f",
        x"0c1fc451fc38",
        x"0c1fc5e1fc51",
        x"0c1fc761fc6a",
        x"0c1fcb51fc83",
        x"0c1fcd31fcc7",
        x"0c200192000b",
        x"0c200262001f",
        x"0c2004520038",
        x"0c2005e20051",
        x"0c200762006a",
        x"0c200b520083",
        x"0c200d3200c7",
        x"0c204192040b",
        x"0c204262041f",
        x"0c2044520438",
        x"0c2045e20451",
        x"0c204762046a",
        x"0c204b520483",
        x"0c204d3204c7",
        x"0c208192080b",
        x"0c2084b2082c",
        x"0c2085720851",
        x"0c208642085e",
        x"0c2088320876",
        x"0c208952088f",
        x"0c208a8208a2",
        x"0c208c1208bb",
        x"0c208d3208c7",
        x"0c20c1920c0b",
        x"0c20c4b20c2c",
        x"0c20c5720c51",
        x"0c20c6420c5e",
        x"0c20c8320c76",
        x"0c20c9520c8f",
        x"0c20ca820ca2",
        x"0c20cc120cbb",
        x"0c20cd320cc7",
        x"0c210192100b",
        x"0c2104b2102c",
        x"0c2105721051",
        x"0c210642105e",
        x"0c2108321076",
        x"0c210952108f",
        x"0c210a8210a2",
        x"0c210c1210bb",
        x"0c210d3210c7",
        x"0c214192140b",
        x"0c2144b2142c",
        x"0c2145721451",
        x"0c214642145e",
        x"0c2148321476",
        x"0c214952148f",
        x"0c214a8214a2",
        x"0c214c1214bb",
        x"0c214d3214c7",
        x"0c218192180b",
        x"0c2184b2182c",
        x"0c2185721851",
        x"0c218642185e",
        x"0c2188321876",
        x"0c218952188f",
        x"0c218a8218a2",
        x"0c218c1218bb",
        x"0c218d3218c7",
        x"0c21c1921c0b",
        x"0c21c4b21c2c",
        x"0c21c5721c51",
        x"0c21c6421c5e",
        x"0c21c8321c76",
        x"0c21c9521c8f",
        x"0c21ca821ca2",
        x"0c21cc121cbb",
        x"0c21cd321cc7",
        x"0c220132200b",
        x"0c2202c22019",
        x"0c220702206a",
        x"0c2207d22076",
        x"0c220ae22089",
        x"0c220c1220bb",
        x"0c220d3220c7",
        x"0c224132240b",
        x"0c2242c22419",
        x"0c224702246a",
        x"0c2247d22476",
        x"0c224ae22489",
        x"0c224c1224bb",
        x"0c224d3224c7",
        x"0c228132280b",
        x"0c2282c22819",
        x"0c228702286a",
        x"0c2287d22876",
        x"0c228ae22889",
        x"0c228c1228bb",
        x"0c228d3228c7",
        x"0c22c1322c0b",
        x"0c22c2c22c19",
        x"0c22c7022c6a",
        x"0c22c7d22c76",
        x"0c22cae22c89",
        x"0c22cc122cbb",
        x"0c22cd322cc7",
        x"0c230132300b",
        x"0c2302c23019",
        x"0c230702306a",
        x"0c2307d23076",
        x"0c230ae23089",
        x"0c230c1230bb",
        x"0c230d3230c7",
        x"0c234132340b",
        x"0c2342c23419",
        x"0c234702346a",
        x"0c2347d23476",
        x"0c234ae23489",
        x"0c234c1234bb",
        x"0c234d3234c7",
        x"0c238192380b",
        x"0c238572384b",
        x"0c2388f23870",
        x"0c2389c23895",
        x"0c238ae238a2",
        x"0c238c1238b5",
        x"0c238d3238c7",
        x"0c23c1923c0b",
        x"0c23c5723c4b",
        x"0c23c8f23c70",
        x"0c23c9c23c95",
        x"0c23cae23ca2",
        x"0c23cc123cb5",
        x"0c23cd323cc7",
        x"0c240192400b",
        x"0c240572404b",
        x"0c2408f24070",
        x"0c2409c24095",
        x"0c240ae240a2",
        x"0c240c1240b5",
        x"0c240d3240c7",
        x"0c244192440b",
        x"0c244572444b",
        x"0c2448f24470",
        x"0c2449c24495",
        x"0c244ae244a2",
        x"0c244c1244b5",
        x"0c244d3244c7",
        x"0c248192480b",
        x"0c248572484b",
        x"0c2488f24870",
        x"0c2489c24895",
        x"0c248ae248a2",
        x"0c248c1248b5",
        x"0c248d3248c7",
        x"0c24c1924c0b",
        x"0c24c5724c4b",
        x"0c24c8f24c70",
        x"0c24c9c24c95",
        x"0c24cae24ca2",
        x"0c24cc124cb5",
        x"0c24cd324cc7",
        x"0c250192500b",
        x"0c250572504b",
        x"0c2508f25070",
        x"0c2509c25095",
        x"0c250ae250a2",
        x"0c250c1250b5",
        x"0c250d3250c7",
        x"0c254192540b",
        x"0c2542c2541f",
        x"0c2544525432",
        x"0c2545e25457",
        x"0c2548325464",
        x"0c254d325495",
        x"0c258192580b",
        x"0c2582c2581f",
        x"0c2584525832",
        x"0c2585e25857",
        x"0c2588325864",
        x"0c258d325895",
        x"0c25c1925c0b",
        x"0c25c2c25c1f",
        x"0c25c4525c32",
        x"0c25c5e25c57",
        x"0c25c8325c64",
        x"0c25cd325c95",
        x"0c260192600b",
        x"0c2602c2601f",
        x"0c2604526032",
        x"0c2605e26057",
        x"0c2608326064",
        x"0c260d326095",
        x"0c264192640b",
        x"0c2642c2641f",
        x"0c2644526432",
        x"0c2645e26457",
        x"0c2648326464",
        x"0c264d326495",
        x"0c268192680b",
        x"0c2682c2681f",
        x"0c2684526832",
        x"0c2685e26857",
        x"0c2688326864",
        x"0c268d326895",
        x"0c26c1f26c0b",
        x"0c26c3826c32",
        x"0c26c4526c3e",
        x"0c26c5726c51",
        x"0c26c6a26c5e",
        x"0c26c8f26c70",
        x"0c26c9c26c95",
        x"0c26cd326cc7",
        x"0c2701f2700b",
        x"0c2703827032",
        x"0c270452703e",
        x"0c2705727051",
        x"0c2706a2705e",
        x"0c2708f27070",
        x"0c2709c27095",
        x"0c270d3270c7",
        x"0c2741f2740b",
        x"0c2743827432",
        x"0c274452743e",
        x"0c2745727451",
        x"0c2746a2745e",
        x"0c2748f27470",
        x"0c2749c27495",
        x"0c274d3274c7",
        x"0c2781f2780b",
        x"0c2783827832",
        x"0c278452783e",
        x"0c2785727851",
        x"0c2786a2785e",
        x"0c2788f27870",
        x"0c2789c27895",
        x"0c278d3278c7",
        x"0c27c1f27c0b",
        x"0c27c3827c32",
        x"0c27c4527c3e",
        x"0c27c5727c51",
        x"0c27c6a27c5e",
        x"0c27c8f27c70",
        x"0c27c9c27c95",
        x"0c27cd327cc7",
        x"0c2801f2800b",
        x"0c2803828032",
        x"0c280452803e",
        x"0c2805728051",
        x"0c2806a2805e",
        x"0c2808f28070",
        x"0c2809c28095",
        x"0c280d3280c7",
        x"0c284132840b",
        x"0c2842c28426",
        x"0c2844528432",
        x"0c284512844b",
        x"0c2846a28457",
        x"0c2847d28476",
        x"0c2849c2848f",
        x"0c284c0284a2",
        x"0c284d3284c7",
        x"0c288132880b",
        x"0c2882c28826",
        x"0c2884528832",
        x"0c288512884b",
        x"0c2886a28857",
        x"0c2887d28876",
        x"0c2889c2888f",
        x"0c288c0288a2",
        x"0c288d3288c7",
        x"0c28c1328c0b",
        x"0c28c2c28c26",
        x"0c28c4528c32",
        x"0c28c5128c4b",
        x"0c28c6a28c57",
        x"0c28c7d28c76",
        x"0c28c9c28c8f",
        x"0c28cc028ca2",
        x"0c28cd328cc7",
        x"0c290132900b",
        x"0c2902c29026",
        x"0c2904529032",
        x"0c290512904b",
        x"0c2906a29057",
        x"0c2907d29076",
        x"0c2909c2908f",
        x"0c290c0290a2",
        x"0c290d3290c7",
        x"0c294132940b",
        x"0c2942c29426",
        x"0c2944529432",
        x"0c294512944b",
        x"0c2946a29457",
        x"0c2947d29476",
        x"0c2949c2948f",
        x"0c294c0294a2",
        x"0c294d3294c7",
        x"0c298132980b",
        x"0c2982c29826",
        x"0c2984529832",
        x"0c298512984b",
        x"0c2986a29857",
        x"0c2987d29876",
        x"0c2989c2988f",
        x"0c298c0298a2",
        x"0c298d3298c7",
        x"0c29c1329c0b",
        x"0c29c2c29c26",
        x"0c29c5129c4b",
        x"0c29c5e29c57",
        x"0c29c8f29c76",
        x"0c29c9c29c95",
        x"0c29ca829ca2",
        x"0c29cc029cbb",
        x"0c29cd329cc7",
        x"0c2a0132a00b",
        x"0c2a02c2a026",
        x"0c2a0512a04b",
        x"0c2a05e2a057",
        x"0c2a08f2a076",
        x"0c2a09c2a095",
        x"0c2a0a82a0a2",
        x"0c2a0c02a0bb",
        x"0c2a0d32a0c7",
        x"0c2a4132a40b",
        x"0c2a42c2a426",
        x"0c2a4512a44b",
        x"0c2a45e2a457",
        x"0c2a48f2a476",
        x"0c2a49c2a495",
        x"0c2a4a82a4a2",
        x"0c2a4c02a4bb",
        x"0c2a4d32a4c7",
        x"0c2a8132a80b",
        x"0c2a82c2a826",
        x"0c2a8512a84b",
        x"0c2a85e2a857",
        x"0c2a88f2a876",
        x"0c2a89c2a895",
        x"0c2a8a82a8a2",
        x"0c2a8c02a8bb",
        x"0c2a8d32a8c7",
        x"0c2ac132ac0b",
        x"0c2ac2c2ac26",
        x"0c2ac512ac4b",
        x"0c2ac5e2ac57",
        x"0c2ac8f2ac76",
        x"0c2ac9c2ac95",
        x"0c2aca82aca2",
        x"0c2acc02acbb",
        x"0c2acd32acc7",
        x"0c2b0132b00b",
        x"0c2b02c2b026",
        x"0c2b0512b04b",
        x"0c2b05e2b057",
        x"0c2b08f2b076",
        x"0c2b09c2b095",
        x"0c2b0a82b0a2",
        x"0c2b0c02b0bb",
        x"0c2b0d32b0c7",
        x"0c2b4322b40b",
        x"0c2b43e2b438",
        x"0c2b45e2b44b",
        x"0c2b47d2b470",
        x"0c2b48f2b483",
        x"0c2b49c2b495",
        x"0c2b4a82b4a2",
        x"0c2b4c02b4bb",
        x"0c2b4d32b4c7",
        x"0c2b8322b80b",
        x"0c2b83e2b838",
        x"0c2b85e2b84b",
        x"0c2b87d2b870",
        x"0c2b88f2b883",
        x"0c2b89c2b895",
        x"0c2b8a82b8a2",
        x"0c2b8c02b8bb",
        x"0c2b8d32b8c7",
        x"0c2bc322bc0b",
        x"0c2bc3e2bc38",
        x"0c2bc5e2bc4b",
        x"0c2bc7d2bc70",
        x"0c2bc8f2bc83",
        x"0c2bc9c2bc95",
        x"0c2bca82bca2",
        x"0c2bcc02bcbb",
        x"0c2bcd32bcc7",
        x"0c2c0322c00b",
        x"0c2c03e2c038",
        x"0c2c05e2c04b",
        x"0c2c07d2c070",
        x"0c2c08f2c083",
        x"0c2c09c2c095",
        x"0c2c0a82c0a2",
        x"0c2c0c02c0bb",
        x"0c2c0d32c0c7",
        x"0c2c4322c40b",
        x"0c2c43e2c438",
        x"0c2c45e2c44b",
        x"0c2c47d2c470",
        x"0c2c48f2c483",
        x"0c2c49c2c495",
        x"0c2c4a82c4a2",
        x"0c2c4c02c4bb",
        x"0c2c4d32c4c7",
        x"0c2c8322c80b",
        x"0c2c83e2c838",
        x"0c2c85e2c84b",
        x"0c2c87d2c870",
        x"0c2c88f2c883",
        x"0c2c89c2c895",
        x"0c2c8a82c8a2",
        x"0c2c8c02c8bb",
        x"0c2c8d32c8c7",
        x"0c2cc322cc0b",
        x"0c2cc3e2cc38",
        x"0c2cc5e2cc4b",
        x"0c2cc7d2cc70",
        x"0c2cc8f2cc83",
        x"0c2cc9c2cc95",
        x"0c2cca82cca2",
        x"0c2ccc02ccbb",
        x"0c2ccd32ccc7",
        x"0c2d0192d00b",
        x"0c2d0322d026",
        x"0c2d04b2d045",
        x"0c2d0572d051",
        x"0c2d0642d05e",
        x"0c2d09c2d095",
        x"0c2d0a82d0a2",
        x"0c2d0c02d0bb",
        x"0c2d0d32d0c7",
        x"0c2d4192d40b",
        x"0c2d4322d426",
        x"0c2d44b2d445",
        x"0c2d4572d451",
        x"0c2d4642d45e",
        x"0c2d49c2d495",
        x"0c2d4a82d4a2",
        x"0c2d4c02d4bb",
        x"0c2d4d32d4c7",
        x"0c2d8192d80b",
        x"0c2d8322d826",
        x"0c2d84b2d845",
        x"0c2d8572d851",
        x"0c2d8642d85e",
        x"0c2d89c2d895",
        x"0c2d8a82d8a2",
        x"0c2d8c02d8bb",
        x"0c2d8d32d8c7",
        x"0c2dc192dc0b",
        x"0c2dc322dc26",
        x"0c2dc4b2dc45",
        x"0c2dc572dc51",
        x"0c2dc642dc5e",
        x"0c2dc9c2dc95",
        x"0c2dca82dca2",
        x"0c2dcc02dcbb",
        x"0c2dcd32dcc7",
        x"0c2e0192e00b",
        x"0c2e0322e026",
        x"0c2e04b2e045",
        x"0c2e0572e051",
        x"0c2e0642e05e",
        x"0c2e09c2e095",
        x"0c2e0a82e0a2",
        x"0c2e0c02e0bb",
        x"0c2e0d32e0c7",
        x"0c2e4192e40b",
        x"0c2e4322e426",
        x"0c2e44b2e445",
        x"0c2e4572e451",
        x"0c2e4642e45e",
        x"0c2e49c2e495",
        x"0c2e4a82e4a2",
        x"0c2e4c02e4bb",
        x"0c2e4d32e4c7",
        x"0c2e8132e80b",
        x"0c2e81f2e819",
        x"0c2e83e2e82c",
        x"0c2e85e2e84b",
        x"0c2e86a2e864",
        x"0c2e87d2e870",
        x"0c2e88f2e889",
        x"0c2e89c2e895",
        x"0c2e8c02e8a2",
        x"0c2e8d32e8c7",
        x"0c2ec132ec0b",
        x"0c2ec1f2ec19",
        x"0c2ec3e2ec2c",
        x"0c2ec5e2ec4b",
        x"0c2ec6a2ec64",
        x"0c2ec7d2ec70",
        x"0c2ec8f2ec89",
        x"0c2ec9c2ec95",
        x"0c2ecc02eca2",
        x"0c2ecd32ecc7",
        x"0c2f0132f00b",
        x"0c2f01f2f019",
        x"0c2f03e2f02c",
        x"0c2f05e2f04b",
        x"0c2f06a2f064",
        x"0c2f07d2f070",
        x"0c2f08f2f089",
        x"0c2f09c2f095",
        x"0c2f0c02f0a2",
        x"0c2f0d32f0c7",
        x"0c2f4132f40b",
        x"0c2f41f2f419",
        x"0c2f43e2f42c",
        x"0c2f45e2f44b",
        x"0c2f46a2f464",
        x"0c2f47d2f470",
        x"0c2f48f2f489",
        x"0c2f49c2f495",
        x"0c2f4c02f4a2",
        x"0c2f4d32f4c7",
        x"0c2f8132f80b",
        x"0c2f81f2f819",
        x"0c2f83e2f82c",
        x"0c2f85e2f84b",
        x"0c2f86a2f864",
        x"0c2f87d2f870",
        x"0c2f88f2f889",
        x"0c2f89c2f895",
        x"0c2f8c02f8a2",
        x"0c2f8d32f8c7",
        x"0c2fc132fc0b",
        x"0c2fc1f2fc19",
        x"0c2fc3e2fc2c",
        x"0c2fc5e2fc4b",
        x"0c2fc6a2fc64",
        x"0c2fc7d2fc70",
        x"0c2fc8f2fc89",
        x"0c2fc9c2fc95",
        x"0c2fcc02fca2",
        x"0c2fcd32fcc7",
        x"0c3001f3000b",
        x"0c3003830032",
        x"0c3005730051",
        x"0c300643005e",
        x"0c300703006a",
        x"0c3008930076",
        x"0c3009c30095",
        x"0c300d3300c7",
        x"0c3041f3040b",
        x"0c3043830432",
        x"0c3045730451",
        x"0c304643045e",
        x"0c304703046a",
        x"0c3048930476",
        x"0c3049c30495",
        x"0c304d3304c7",
        x"0c3081f3080b",
        x"0c3083830832",
        x"0c3085730851",
        x"0c308643085e",
        x"0c308703086a",
        x"0c3088930876",
        x"0c3089c30895",
        x"0c308d3308c7",
        x"0c30c1f30c0b",
        x"0c30c3830c32",
        x"0c30c5730c51",
        x"0c30c6430c5e",
        x"0c30c7030c6a",
        x"0c30c8930c76",
        x"0c30c9c30c95",
        x"0c30cd330cc7",
        x"0c3101f3100b",
        x"0c3103831032",
        x"0c3105731051",
        x"0c310643105e",
        x"0c310703106a",
        x"0c3108931076",
        x"0c3109c31095",
        x"0c310d3310c7",
        x"0c3141f3140b",
        x"0c3143831432",
        x"0c3145731451",
        x"0c314643145e",
        x"0c314703146a",
        x"0c3148931476",
        x"0c3149c31495",
        x"0c314d3314c7",
        x"0c318d33180b",
        x"0c31cd331c0b",
        x"0c320d33200b",
        x"0c324d33240b",                --fin qr
        OTHERS => x"000000000000");
BEGIN

    PROCESS(clk)
    BEGIN
        IF falling_edge(clk) THEN
            IF ce = '1' THEN
                data_out_read_only <= memory_data(to_integer(unsigned(address_read_only)));
                IF rw = '1' THEN        -- write
                    memory_data(to_integer(unsigned(address))) <= input;
                ELSE                    --read
                    data_out <= memory_data(to_integer(unsigned(address)));
                END IF;
            END IF;
        END IF;
    END PROCESS;

END Behavioral;
