----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08.02.2023 15:29:34
-- Design Name: 
-- Module Name: graphic_memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY graphic_memory IS
    PORT(
        clk                : IN  STD_LOGIC;
        ce                 : IN  STD_LOGIC;
        rw                 : IN  STD_LOGIC; --R/=0 W=1
        address_read_only  : IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
        address            : IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
        input              : IN  STD_LOGIC_VECTOR(47 DOWNTO 0);
        data_out_read_only : OUT STD_LOGIC_VECTOR(47 DOWNTO 0);
        data_out           : OUT STD_LOGIC_VECTOR(47 DOWNTO 0));
END graphic_memory;

ARCHITECTURE Behavioral OF graphic_memory IS
    TYPE memory_array IS ARRAY (INTEGER RANGE 0 TO 4095) OF STD_LOGIC_VECTOR(47 DOWNTO 0);
    SIGNAL memory_data : memory_array := ( --x/y
    x"0c4c4094c407",--debut graph
x"0c4c40f4c40b",
x"0c4c4134c411",
x"0c4c8094c806",
x"0c4c80f4c80b",
x"0c4c8144c810",
x"0c4cc084cc06",
x"0c4cc0d4cc0b",
x"0c4cc114cc10",
x"0c4cc154cc13",
x"0c4ce6d4cc17",
x"0c4d00a4d006",
x"0c4d00f4d00b",
x"0c4d0114d010",
x"0c4d0154d013",
x"0c4d26d4d017",
x"0c4d4074d406",
x"0c4d40a4d409",
x"0c4d40f4d40d",
x"0c4d4114d410",
x"0c4d4154d413",
x"0c4d66d4d417",
x"0c4d80a4d806",
x"0c4d80c4d80b",
x"0c4d80f4d80d",
x"0c4d8144d810",
x"0c4d8194d817",
x"0c4d87d4d87a",
x"0c4d8e04d8dd",
x"0c4d9434d941",
x"0c4d9a74d9a4",
x"0c4da0a4da07",
x"0c4da6d4da6a",
x"0c4dc094dc06",
x"0c4dc0e4dc0b",
x"0c4dc144dc11",
x"0c4dc194dc17",
x"0c4dc7d4dc7a",
x"0c4dce04dcdd",
x"0c4dd434dd41",
x"0c4dda74dda4",
x"0c4de0a4de07",
x"0c4de6d4de6a",
x"0c4e0194e017",
x"0c4e07d4e07a",
x"0c4e0e04e0dd",
x"0c4e1434e141",
x"0c4e1a74e1a4",
x"0c4e20a4e207",
x"0c4e26d4e26a",
x"0c4e4194e417",
x"0c4e47d4e47a",
x"0c4e4e04e4dd",
x"0c4e5434e541",
x"0c4e5a74e5a4",
x"0c4e60a4e607",
x"0c4e66d4e66a",
x"0c4e8194e817",
x"0c4e87d4e87a",
x"0c4e8e04e8dd",
x"0c4e9434e941",
x"0c4e9a74e9a4",
x"0c4ea0a4ea07",
x"0c4ea6d4ea6a",
x"0c4ec194ec17",
x"0c4ee6d4ee6a",
x"0c4f0194f017",
x"0c4f26d4f26a",
x"0c4f4194f417",
x"0c4f66d4f66a",
x"0c4f8194f817",
x"0c4fa6d4fa6a",
x"0c4fc194fc17",
x"0c4fe6d4fe6a",
x"0c5001950017",
x"0c5026d5026a",
x"0c5041950417",
x"0c5066d5066a",
x"0c5081950817",
x"0c50a6d50a6a",
x"0c50c1950c17",
x"0c50e6d50e6a",
x"0c5101951017",
x"0c5126951259",
x"0c5126d5126a",
x"0c5141951417",
x"0c5166951658",
x"0c5166d5166a",
x"0c5181951817",
x"0c51a6951a57",
x"0c51a6d51a6a",
x"0c51c1951c17",
x"0c51e5a51e57",
x"0c51e6d51e6a",
x"0c5201952017",
x"0c5225952256",
x"0c5226d5226a",
x"0c5241952417",
x"0c5265952655",
x"0c5266d5266a",
x"0c5281952817",
x"0c52a5852a55",
x"0c52a6d52a6a",
x"0c52c1952c17",
x"0c52e5852e54",
x"0c52e6d52e6a",
x"0c5301953017",
x"0c5325753235",
x"0c5326d5326a",
x"0c5341953417",
x"0c5365653634",
x"0c5366d5366a",
x"0c5381953817",
x"0c53a5653a34",
x"0c53a6d53a6a",
x"0c53c1953c17",
x"0c53e3753e34",
x"0c53e6d53e6a",
x"0c5401954017",
x"0c5423754233",
x"0c5426d5426a",
x"0c5441954417",
x"0c5463654633",
x"0c5466d5466a",
x"0c5480b54807",
x"0c548105480c",
x"0c5481554811",
x"0c5481954817",
x"0c54a3654a33",
x"0c54a6d54a6a",
x"0c54c0854c07",
x"0c54c0d54c0c",
x"0c54c1254c0e",
x"0c54c1554c13",
x"0c54c1954c17",
x"0c54e3654e33",
x"0c54e6d54e6a",
x"0c5500d55007",
x"0c550125500f",
x"0c5501555014",
x"0c5501e55017",
x"0c5523655217",
x"0c5526d55265",
x"0c5540d55407",
x"0c554125540f",
x"0c5541555414",
x"0c5541f55417",
x"0c5563555616",
x"0c5566d55665",
x"0c5580855807",
x"0c5580d55809",
x"0c558125580e",
x"0c5581555813",
x"0c5581e55817",
x"0c55a3555a16",
x"0c55a6d55a65",
x"0c55c0b55c07",
x"0c55c1055c0c",
x"0c55c1555c11",
x"0c55c1955c17",
x"0c55e1955e15",
x"0c55e6d55e6a",
x"0c5600956008",
x"0c5600f5600d",
x"0c5601456012",
x"0c5601956017",
x"0c5621856214",
x"0c5626d5626a",
x"0c5641956417",
x"0c5661756614",
x"0c5666d5666a",
x"0c5681956817",
x"0c56a1756a13",
x"0c56a6d56a6a",
x"0c56c1956c17",
x"0c56e1656e13",
x"0c56e6d56e6a",
x"0c5701957017",
x"0c57216571f8",
x"0c5726d5726a",
x"0c5741957417",
x"0c57615575f7",
x"0c5766d5766a",
x"0c5781957817",
x"0c57a14579f6",
x"0c57a6d57a6a",
x"0c57c1957c17",
x"0c57dfa57df6",
x"0c57e6d57e6a",
x"0c5801958017",
x"0c581f9581f5",
x"0c5826d5826a",
x"0c5841958417",
x"0c585f8585f5",
x"0c5866d5866a",
x"0c5881958817",
x"0c589f8589f5",
x"0c58a6d58a6a",
x"0c58c1958c17",
x"0c58df858df4",
x"0c58e6d58e6a",
x"0c5901959017",
x"0c591f7591da",
x"0c5926d5926a",
x"0c5941959417",
x"0c595f7595d9",
x"0c5966d5966a",
x"0c5981959817",
x"0c599f6599d7",
x"0c59a6d59a6a",
x"0c59c1959c17",
x"0c59ddb59dd6",
x"0c59e6d59e6a",
x"0c5a0195a017",
x"0c5a1da5a1d5",
x"0c5a26d5a26a",
x"0c5a4195a417",
x"0c5a5d85a5d4",
x"0c5a66d5a66a",
x"0c5a8195a817",
x"0c5a9d75a9d2",
x"0c5aa6d5aa6a",
x"0c5ac195ac17",
x"0c5add65add1",
x"0c5ae6d5ae6a",
x"0c5b0195b017",
x"0c5b1d55b1bf",
x"0c5b26d5b26a",
x"0c5b4195b417",
x"0c5b5d35b5be",
x"0c5b66d5b66a",
x"0c5b8195b817",
x"0c5b9d25b9bd",
x"0c5ba6d5ba6a",
x"0c5bc195bc17",
x"0c5bdc15bdbd",
x"0c5be6d5be6a",
x"0c5c0195c017",
x"0c5c1c05c1bc",
x"0c5c26d5c26a",
x"0c5c4195c417",
x"0c5c5bf5c5bb",
x"0c5c66d5c66a",
x"0c5c8195c817",
x"0c5c9be5c9ba",
x"0c5ca6d5ca6a",
x"0c5cc195cc17",
x"0c5cdbd5cdb9",
x"0c5ce6d5ce6a",
x"0c5d0095d005",
x"0c5d00f5d00b",
x"0c5d0135d010",
x"0c5d0195d017",
x"0c5d1bd5d1b9",
x"0c5d26d5d26a",
x"0c5d4075d405",
x"0c5d40c5d40b",
x"0c5d4115d40f",
x"0c5d4145d412",
x"0c5d41a5d417",
x"0c5d5bc5d59d",
x"0c5d66d5d66a",
x"0c5d8095d805",
x"0c5d80e5d80b",
x"0c5d8115d80f",
x"0c5d8145d813",
x"0c5d81f5d817",
x"0c5d9bb5d99c",
x"0c5da6d5da65",
x"0c5dc0a5dc07",
x"0c5dc115dc0c",
x"0c5dc145dc13",
x"0c5dc1f5dc17",
x"0c5dda05dd9b",
x"0c5ddba5ddb9",
x"0c5de6d5de65",
x"0c5e00a5e008",
x"0c5e0115e00d",
x"0c5e0145e012",
x"0c5e01e5e017",
x"0c5e19f5e19b",
x"0c5e26d5e265",
x"0c5e4095e405",
x"0c5e40e5e40a",
x"0c5e4145e410",
x"0c5e4195e417",
x"0c5e59e5e59a",
x"0c5e66d5e66a",
x"0c5e8085e806",
x"0c5e80d5e80b",
x"0c5e8135e811",
x"0c5e8195e817",
x"0c5e99d5e999",
x"0c5ea6d5ea6a",
x"0c5ec195ec17",
x"0c5ed9c5ed98",
x"0c5ee6d5ee6a",
x"0c5f0195f017",
x"0c5f19b5f197",
x"0c5f26d5f26a",
x"0c5f4195f417",
x"0c5f59a5f583",
x"0c5f66d5f66a",
x"0c5f8195f817",
x"0c5f99a5f982",
x"0c5fa6d5fa6a",
x"0c5fc195fc17",
x"0c5fd865fd82",
x"0c5fd985fd87",
x"0c5fe6d5fe6a",
x"0c6001960017",
x"0c6018560181",
x"0c6026d6026a",
x"0c6041960417",
x"0c6058460581",
x"0c6066d6066a",
x"0c6081960817",
x"0c6098460981",
x"0c60a6d60a6a",
x"0c60c1960c17",
x"0c60d8460d80",
x"0c60e6d60e6a",
x"0c6101961017",
x"0c6118361180",
x"0c6126d6126a",
x"0c6141961417",
x"0c6158361567",
x"0c6166d6166a",
x"0c6181961817",
x"0c6198261966",
x"0c61a6d61a6a",
x"0c61c1961c17",
x"0c61d6a61d66",
x"0c61d8161d6b",
x"0c61e6d61e6a",
x"0c6201962017",
x"0c6216962166",
x"0c6226d6226a",
x"0c6241962417",
x"0c6256962566",
x"0c6266d6266a",
x"0c6281962817",
x"0c6296962965",
x"0c62a6d62a6a",
x"0c62c1962c17",
x"0c62d6862d65",
x"0c62e6d62e6a",
x"0c6301963017",
x"0c6316863165",
x"0c6326d6326a",
x"0c6341963417",
x"0c6356863550",
x"0c6366d6366a",
x"0c6381963817",
x"0c639686394f",
x"0c63a6d63a6a",
x"0c63c1963c17",
x"0c63d6763d4e",
x"0c63e6d63e6a",
x"0c6401964017",
x"0c641516414e",
x"0c6426d6426a",
x"0c6441964417",
x"0c645516454d",
x"0c6466d6466a",
x"0c6481964817",
x"0c649506494c",
x"0c64a6d64a6a",
x"0c64c1964c17",
x"0c64d4f64d4b",
x"0c64e6d64e6a",
x"0c6501965017",
x"0c6514f6514b",
x"0c6526d6526a",
x"0c6540b65407",
x"0c654106540d",
x"0c6541565412",
x"0c6541965417",
x"0c6554e65535",
x"0c6566d6566a",
x"0c6580965807",
x"0c6580e6580c",
x"0c658136580f",
x"0c6581565814",
x"0c6581965817",
x"0c6594d65935",
x"0c65a6d65a6a",
x"0c65c0965c07",
x"0c65c0d65c0c",
x"0c65c1365c0f",
x"0c65c1665c14",
x"0c65c1a65c17",
x"0c65d4c65d34",
x"0c65e6d65e6a",
x"0c6600b66007",
x"0c6600d6600c",
x"0c660136600f",
x"0c6601666014",
x"0c6601f66017",
x"0c6613766134",
x"0c6626d66265",
x"0c6640d6640a",
x"0c664136640f",
x"0c6641666414",
x"0c6641f66417",
x"0c6653766533",
x"0c6666d66665",
x"0c6680b66807",
x"0c668106680c",
x"0c6681566811",
x"0c6681a66817",
x"0c6693766933",
x"0c66a6d66a6a",
x"0c66c0a66c07",
x"0c66c0f66c0d",
x"0c66c1466c12",
x"0c66c1966c17",
x"0c66d3666d33",
x"0c66e6d66e6a",
x"0c6701967017",
x"0c6713667132",
x"0c6726d6726a",
x"0c6741967417",
x"0c6753567524",
x"0c6766d6766a",
x"0c6781967817",
x"0c6793567923",
x"0c67a6d67a6a",
x"0c67c1967c17",
x"0c67d3467d22",
x"0c67e6d67e6a",
x"0c6801968017",
x"0c6812568121",
x"0c6826d6826a",
x"0c6841968417",
x"0c6852468520",
x"0c6866d6866a",
x"0c6881968817",
x"0c6892368920",
x"0c68a6d68a6a",
x"0c68c1968c17",
x"0c68d2368d1f",
x"0c68e6d68e6a",
x"0c6901969017",
x"0c691226911e",
x"0c6926d6926a",
x"0c6941969417",
x"0c6952169509",
x"0c6966d6966a",
x"0c6981969817",
x"0c6992069908",
x"0c69a6d69a6a",
x"0c69c1969c17",
x"0c69d1f69d07",
x"0c69e6d69e6a",
x"0c6a0196a017",
x"0c6a10a6a107",
x"0c6a26d6a26a",
x"0c6a4196a417",
x"0c6a50a6a506",
x"0c6a66d6a66a",
x"0c6a8196a817",
x"0c6a9096a906",
x"0c6aa6d6aa6a",
x"0c6ac196ac17",
x"0c6ad096ad05",
x"0c6ae6d6ae6a",
x"0c6b0196b017",
x"0c6b1086b105",
x"0c6b26d6b26a",
x"0c6b4196b417",
x"0c6b5086b4f3",
x"0c6b66d6b66a",
x"0c6b8196b817",
x"0c6b9076b8f2",
x"0c6ba6d6ba6a",
x"0c6bc196bc17",
x"0c6bd076bcf2",
x"0c6be6d6be6a",
x"0c6c0196c017",
x"0c6c0f56c0f2",
x"0c6c26d6c26a",
x"0c6c4196c417",
x"0c6c4f56c4f1",
x"0c6c66d6c66a",
x"0c6c8196c817",
x"0c6c8f56c8f1",
x"0c6ca6d6ca6a",
x"0c6cc196cc17",
x"0c6ccf46ccf1",
x"0c6ce6d6ce6a",
x"0c6d0196d017",
x"0c6d0f46d0f1",
x"0c6d26d6d26a",
x"0c6d4196d417",
x"0c6d4f46d4de",
x"0c6d66d6d66a",
x"0c6d8196d817",
x"0c6d8f36d8dd",
x"0c6da6d6da6a",
x"0c6dc0b6dc09",
x"0c6dc116dc0d",
x"0c6dc156dc12",
x"0c6dc196dc17",
x"0c6dcf36dcdd",
x"0c6de6d6de6a",
x"0c6e00b6e009",
x"0c6e00e6e00d",
x"0c6e0166e012",
x"0c6e0196e017",
x"0c6e0e06e0dd",
x"0c6e26d6e26a",
x"0c6e40b6e408",
x"0c6e40f6e40d",
x"0c6e4136e411",
x"0c6e41e6e414",
x"0c6e4e06e4dd",
x"0c6e66d6e665",
x"0c6e8096e807",
x"0c6e80b6e80a",
x"0c6e8106e80d",
x"0c6e8136e811",
x"0c6e81f6e815",
x"0c6e8e06e8dc",
x"0c6ea6d6ea65",
x"0c6ec0c6ec07",
x"0c6ec136ec0f",
x"0c6ec1e6ec14",
x"0c6ecdf6ecdc",
x"0c6ee6d6ee65",
x"0c6f0116f009",
x"0c6f0166f012",
x"0c6f0196f017",
x"0c6f0df6f0dc",
x"0c6f26d6f26a",
x"0c6f40b6f40a",
x"0c6f4106f40d",
x"0c6f4156f412",
x"0c6f4196f417",
x"0c6f4df6f4cd",
x"0c6f66d6f66a",
x"0c6f8196f817",
x"0c6f8df6f8cc",
x"0c6fa6d6fa6a",
x"0c6fc196fc17",
x"0c6fcde6fccc",
x"0c6fe6d6fe6a",
x"0c7001970017",
x"0c700cf700cc",
x"0c7026d7026a",
x"0c7041970417",
x"0c704cf704cb",
x"0c7066d7066a",
x"0c7081970817",
x"0c708ce708cb",
x"0c70a6d70a6a",
x"0c70c1970c17",
x"0c70cce70ccb",
x"0c70e6d70e6a",
x"0c7101971017",
x"0c710ce710ca",
x"0c7126d7126a",
x"0c7141971417",
x"0c714cd714bc",
x"0c7166d7166a",
x"0c7181971817",
x"0c718cd718bb",
x"0c71a6d71a6a",
x"0c71c1971c17",
x"0c71ccc71cba",
x"0c71e6d71e6a",
x"0c7201972017",
x"0c720bd720b9",
x"0c7226d7226a",
x"0c7241972417",
x"0c724bc724b8",
x"0c7266d7266a",
x"0c7281972817",
x"0c728bb728b7",
x"0c72a6d72a6a",
x"0c72c1972c17",
x"0c72cba72cb6",
x"0c72e6d72e6a",
x"0c7301973017",
x"0c730b9730b5",
x"0c7326d7326a",
x"0c7341973417",
x"0c734b8734a9",
x"0c7366d7366a",
x"0c7381973817",
x"0c738b7738a8",
x"0c73a6d73a6a",
x"0c73c1973c17",
x"0c73cb773ca8",
x"0c73e6d73e6a",
x"0c7401974017",
x"0c740ab740a7",
x"0c7426d7426a",
x"0c7441974417",
x"0c744aa744a7",
x"0c7466d7466a",
x"0c7481974817",
x"0c748aa748a7",
x"0c74a6d74a6a",
x"0c74c1974c17",
x"0c74caa74ca6",
x"0c74e6d74e6a",
x"0c7501975017",
x"0c750aa750a6",
x"0c7526d7526a",
x"0c7541975417",
x"0c754a975497",
x"0c7566d7566a",
x"0c7581975817",
x"0c758a975896",
x"0c75a6d75a6a",
x"0c75c1975c17",
x"0c75ca975c96",
x"0c75e6d75e6a",
x"0c7600b76009",
x"0c760107600d",
x"0c7601476012",
x"0c7601976017",
x"0c7609976095",
x"0c7626d7626a",
x"0c7640b76408",
x"0c764107640c",
x"0c7641576411",
x"0c7641976417",
x"0c7649876495",
x"0c7666d7666a",
x"0c7680b76808",
x"0c7680d7680c",
x"0c768137680f",
x"0c7681676814",
x"0c7681a76817",
x"0c7689876894",
x"0c76a6d76a6a",
x"0c76c0b76c07",
x"0c76c0d76c0c",
x"0c76c1376c0f",
x"0c76c1676c14",
x"0c76c1f76c17",
x"0c76c9776c94",
x"0c76e6d76e65",
x"0c7700d77007",
x"0c770137700f",
x"0c7701677014",
x"0c7701f77017",
x"0c7709777094",
x"0c7726d77265",
x"0c7741077407",
x"0c7741377411",
x"0c7741577414",
x"0c7741e77417",
x"0c7749777488",
x"0c7766d77666",
x"0c7780b77809",
x"0c778107780d",
x"0c7781577812",
x"0c7781977817",
x"0c7789677887",
x"0c77a6d77a6a",
x"0c77c1977c17",
x"0c77c9677c87",
x"0c77e6d77e6a",
x"0c7801978017",
x"0c7808a78087",
x"0c7826d7826a",
x"0c7841978417",
x"0c7848a78486",
x"0c7866d7866a",
x"0c7881978817",
x"0c7888978886",
x"0c78a6d78a6a",
x"0c78c1978c17",
x"0c78c8978c86",
x"0c78e6d78e6a",
x"0c7901979017",
x"0c7908979086",
x"0c7926d7926a",
x"0c7941979417",
x"0c7948879479",
x"0c7966d7966a",
x"0c7981979817",
x"0c7988879878",
x"0c79a6d79a6a",
x"0c79c1979c17",
x"0c79c8879c78",
x"0c79e6d79e6a",
x"0c7a0197a017",
x"0c7a07b7a078",
x"0c7a26d7a26a",
x"0c7a4197a417",
x"0c7a47b7a477",
x"0c7a66d7a66a",
x"0c7a8197a817",
x"0c7a87a7a877",
x"0c7aa6d7aa6a",
x"0c7ac197ac17",
x"0c7ac7a7ac77",
x"0c7ae6d7ae6a",
x"0c7b0197b017",
x"0c7b07a7b077",
x"0c7b26d7b26a",
x"0c7b4197b417",
x"0c7b47a7b476",
x"0c7b66d7b66a",
x"0c7b8197b817",
x"0c7b8797b86c",
x"0c7ba6d7ba6a",
x"0c7bc197bc17",
x"0c7bc797bc6c",
x"0c7be6d7be6a",
x"0c7c0197c017",
x"0c7c0707c06c",
x"0c7c26d7c26a",
x"0c7c4197c417",
x"0c7c46f7c46c",
x"0c7c66d7c66a",
x"0c7c8197c817",
x"0c7c86f7c86b",
x"0c7ca6d7ca6a",
x"0c7cc197cc17",
x"0c7cc6e7cc6b",
x"0c7ce6d7ce6a",
x"0c7d0197d017",
x"0c7d06e7d06b",
x"0c7d26d7d26a",
x"0c7d4197d417",
x"0c7d46e7d46a",
x"0c7d66d7d66a",
x"0c7d8197d817",
x"0c7d86e7d860",
x"0c7da6d7da6a",
x"0c7dc197dc17",
x"0c7dc6d7dc60",
x"0c7de6d7de6a",
x"0c7e0197e017",
x"0c7e0637e05f",
x"0c7e26d7e26a",
x"0c7e4197e417",
x"0c7e4627e45f",
x"0c7e66d7e66a",
x"0c7e8197e817",
x"0c7e8617e85e",
x"0c7ea6d7ea6a",
x"0c7ec0b7ec07",
x"0c7ec117ec0d",
x"0c7ec157ec12",
x"0c7ec197ec17",
x"0c7ec617ec5d",
x"0c7ee6d7ee6a",
x"0c7f00b7f00a",
x"0c7f00e7f00d",
x"0c7f0137f011",
x"0c7f0167f014",
x"0c7f01e7f017",
x"0c7f0607f05d",
x"0c7f26d7f266",
x"0c7f40b7f408",
x"0c7f4107f40d",
x"0c7f4137f411",
x"0c7f41f7f415",
x"0c7f4607f45c",
x"0c7f66d7f665",
x"0c7f80c7f808",
x"0c7f8137f80e",
x"0c7f81f7f815",
x"0c7f85f7f856",
x"0c7fa6d7fa65",
x"0c7fc0c7fc0a",
x"0c7fc137fc0f",
x"0c7fc1a7fc14",
x"0c7fc5e7fc55",
x"0c7fe6d7fe6a",
x"0c8001080007",
x"0c8001680012",
x"0c8001980017",
x"0c8005880055",
x"0c8026d8026a",
x"0c8040a80408",
x"0c8040f8040d",
x"0c8041580413",
x"0c8041980417",
x"0c8045880454",
x"0c8066d8066a",
x"0c8081980817",
x"0c8085780854",
x"0c80a6d80a6a",
x"0c80c1980c17",
x"0c80c5780c54",
x"0c80e6d80e6a",
x"0c8101981017",
x"0c8105781053",
x"0c8126d8126a",
x"0c8141981417",
x"0c8145681453",
x"0c8166d8166a",
x"0c8181981817",
x"0c8185681849",
x"0c81a6d81a6a",
x"0c81c1981c17",
x"0c81c5581c48",
x"0c81e6d81e6a",
x"0c8201982017",
x"0c8205482048",
x"0c8226d8226a",
x"0c8241982417",
x"0c8244b82448",
x"0c8266d8266a",
x"0c8281982817",
x"0c8284b82848",
x"0c82a6d82a6a",
x"0c82c1982c17",
x"0c82c4b82c47",
x"0c82e6d82e6a",
x"0c8301983017",
x"0c8304a83047",
x"0c8326d8326a",
x"0c8341983417",
x"0c8344a83447",
x"0c8366d8366a",
x"0c8381983817",
x"0c8384a83840",
x"0c83a6d83a6a",
x"0c83c1983c17",
x"0c83c4983c3f",
x"0c83e6d83e6a",
x"0c8401984017",
x"0c840498403f",
x"0c8426d8426a",
x"0c8441984417",
x"0c844428443f",
x"0c8466d8466a",
x"0c8481984817",
x"0c848428483f",
x"0c84a6d84a6a",
x"0c84c1984c17",
x"0c84c4284c3e",
x"0c84e6d84e6a",
x"0c8501985017",
x"0c850418503e",
x"0c8526d8526a",
x"0c8541985417",
x"0c854418543e",
x"0c8566d8566a",
x"0c8581985817",
x"0c8584185838",
x"0c85a6d85a6a",
x"0c85c1985c17",
x"0c85c4185c37",
x"0c85e6d85e6a",
x"0c8601986017",
x"0c8604086037",
x"0c8626d8626a",
x"0c8641986417",
x"0c8643a86437",
x"0c8666d8666a",
x"0c8681986817",
x"0c8683a86836",
x"0c86a6d86a6a",
x"0c86c0a86c07",
x"0c86c0f86c0d",
x"0c86c1486c12",
x"0c86c1986c17",
x"0c86c3986c36",
x"0c86e6d86e6a",
x"0c8700887007",
x"0c8700b87009",
x"0c870108700c",
x"0c8701587011",
x"0c8701987017",
x"0c8703987036",
x"0c8726d8726a",
x"0c8740d87409",
x"0c874128740f",
x"0c8741587414",
x"0c8741987417",
x"0c8743987435",
x"0c8766d8766a",
x"0c8780a87807",
x"0c8780d8780b",
x"0c878128780f",
x"0c8781587814",
x"0c8781e87817",
x"0c8783887831",
x"0c87a6d87a65",
x"0c87c0d87c09",
x"0c87c1287c0f",
x"0c87c1587c14",
x"0c87c1f87c17",
x"0c87c3887c31",
x"0c87e6d87e65",
x"0c8800888007",
x"0c8800b88009",
x"0c880108800c",
x"0c8801588011",
x"0c8801e88017",
x"0c8803788030",
x"0c8826d88265",
x"0c8840a88407",
x"0c8840f8840c",
x"0c8841488411",
x"0c8841988417",
x"0c8843388430",
x"0c8866d8866a",
x"0c8881988817",
x"0c8883388830",
x"0c88a6d88a6a",
x"0c88c1988c17",
x"0c88c3388c2f",
x"0c88e6d88e6a",
x"0c8901989017",
x"0c890328902f",
x"0c8926d8926a",
x"0c8941989417",
x"0c894328942f",
x"0c8966d8966a",
x"0c8981989817",
x"0c8983289829",
x"0c89a6d89a6a",
x"0c89c1989c17",
x"0c89c3289c29",
x"0c89e6d89e6a",
x"0c8a0198a017",
x"0c8a0318a028",
x"0c8a26d8a26a",
x"0c8a4198a417",
x"0c8a42b8a428",
x"0c8a66d8a66a",
x"0c8a8198a817",
x"0c8a82b8a827",
x"0c8aa6d8aa6a",
x"0c8ac198ac17",
x"0c8ac2a8ac27",
x"0c8ae6d8ae6a",
x"0c8b0198b017",
x"0c8b02a8b027",
x"0c8b26d8b26a",
x"0c8b4198b417",
x"0c8b42a8b426",
x"0c8b66d8b66a",
x"0c8b8198b817",
x"0c8b8298b825",
x"0c8ba6d8ba6a",
x"0c8bc198bc17",
x"0c8bc298bc25",
x"0c8be6d8be6a",
x"0c8c0198c017",
x"0c8c0288c024",
x"0c8c26d8c26a",
x"0c8c4198c417",
x"0c8c4278c424",
x"0c8c66d8c66a",
x"0c8c8198c817",
x"0c8c8278c824",
x"0c8ca6d8ca6a",
x"0c8cc198cc17",
x"0c8cc278cc24",
x"0c8ce6d8ce6a",
x"0c8d0198d017",
x"0c8d0278d023",
x"0c8d26d8d26a",
x"0c8d4198d417",
x"0c8d4268d423",
x"0c8d66d8d66a",
x"0c8d8198d817",
x"0c8d8268d81f",
x"0c8da6d8da6a",
x"0c8dc198dc17",
x"0c8dc268dc1f",
x"0c8de6d8de6a",
x"0c8e0198e017",
x"0c8e0258e01e",
x"0c8e26d8e26a",
x"0c8e4198e417",
x"0c8e4218e41e",
x"0c8e66d8e66a",
x"0c8e8198e817",
x"0c8e8218e81e",
x"0c8ea6d8ea6a",
x"0c8ec198ec17",
x"0c8ec218ec1e",
x"0c8ee6d8ee6a",
x"0c8f0198f017",
x"0c8f0218f01d",
x"0c8f26d8f26a",
x"0c8f4198f417",
x"0c8f4208f41d",
x"0c8f66d8f66a",
x"0c8f80a8f807",
x"0c8f8108f80c",
x"0c8f8148f811",
x"0c8f8198f817",
x"0c8f8208f81c",
x"0c8fa6d8fa6a",
x"0c8fc0b8fc07",
x"0c8fc0e8fc0c",
x"0c8fc158fc11",
x"0c8fc1a8fc17",
x"0c8fc208fc1c",
x"0c8fe6d8fe6a",
x"0c9000b90009",
x"0c9000e9000c",
x"0c9001290011",
x"0c9001590014",
x"0c9001f90017",
x"0c9026d90265",
x"0c9040a90408",
x"0c904109040c",
x"0c9041290411",
x"0c9041590414",
x"0c9041f90417",
x"0c9066d90665",
x"0c9080990807",
x"0c908129080e",
x"0c9081590814",
x"0c9081f90817",
x"0c90a6d90a66",
x"0c90c1090c07",
x"0c90c1590c11",
x"0c90c1990c17",
x"0c90c1e90c1b",
x"0c90e6d90e6a",
x"0c9100b91007",
x"0c9100f9100c",
x"0c9101491012",
x"0c9101991017",
x"0c9101e9101b",
x"0c9126d9126a",
x"0c9141991417",
x"0c9141e9141b",
x"0c9166d9166a",
x"0c9181e91817",
x"0c91a6d91a6a",
x"0c91c1e91c17",
x"0c91e6d91e6a",
x"0c9201d92017",
x"0c9226d9226a",
x"0c9241c92417",
x"0c9266d9266a",
x"0c9281c92817",
x"0c92a6d92a6a",
x"0c92c1c92c17",
x"0c92e6d92e6a",
x"0c9301b93017",
x"0c9326d9326a",
x"0c9341b93417",
x"0c9366d9366a",
x"0c9381b93817",
x"0c93a6d93a6a",
x"0c93c1b93c17",
x"0c93e6d93e6a",
x"0c9401b94017",
x"0c9426d9426a",
x"0c9441a94417",
x"0c9466d9466a",
x"0c9481994817",
x"0c94a6d94a6a",
x"0c94c1994c17",
x"0c94e6d94e6a",
x"0c9501995017",
x"0c9526d9526a",
x"0c9541995417",
x"0c9566d9566a",
x"0c9581995817",
x"0c95a6d95a6a",
x"0c95c1995c17",
x"0c95e6d95e6a",
x"0c9601996017",
x"0c9626d9626a",
x"0c9641996417",
x"0c9666d9666a",
x"0c9681996817",
x"0c96a6d96a6a",
x"0c96c1996c17",
x"0c96e6d96e6a",
x"0c9701997017",
x"0c9707d9707a",
x"0c970e0970dd",
x"0c9714397141",
x"0c971a7971a4",
x"0c9720a97207",
x"0c9726d9726a",
x"0c9741997417",
x"0c9747d9747a",
x"0c974e0974dd",
x"0c9754397541",
x"0c975a7975a4",
x"0c9760a97607",
x"0c9766d9766a",
x"0c9780a97806",
x"0c9780f9780b",
x"0c9781497810",
x"0c9781997817",
x"0c9787d9787a",
x"0c978e0978dd",
x"0c9794397941",
x"0c979a7979a4",
x"0c97a0a97a07",
x"0c97a6d97a6a",
x"0c97c0a97c08",
x"0c97c0c97c0b",
x"0c97c1297c0e",
x"0c97c1497c13",
x"0c97c1997c17",
x"0c97c7d97c7a",
x"0c97ce097cdd",
x"0c97d4397d41",
x"0c97da797da4",
x"0c97e0a97e07",
x"0c97e6d97e6a",
x"0c9800a98008",
x"0c9800c9800b",
x"0c980119800e",
x"0c9801598013",
x"0c9801998017",
x"0c9807d9807a",
x"0c980e0980dd",
x"0c9814398141",
x"0c981a7981a4",
x"0c9820a98207",
x"0c9826d9826a",
x"0c9840998407",
x"0c9840c9840b",
x"0c984119840e",
x"0c9841598413",
x"0c9866d98417",
x"0c9880898806",
x"0c9880c9880b",
x"0c9880f9880e",
x"0c9881198810",
x"0c9881498813",
x"0c98a6d98817",
x"0c98c0a98c06",
x"0c98c0f98c0b",
x"0c98c1498c10",
x"0c98e6d98c17",
x"0c9900a99006",
x"0c9900e9900c",
x"0c9901399011",
x"0c9960599603",
x"0c9960a99608",
x"0c9960f9960d",
x"0c9961499612",
x"0c9966399662",
x"0c9966899666",
x"0c9966e9966b",
x"0c9967399670",
x"0c9981a99816",
x"0c9987899875",
x"0c9987d9987a",
x"0c998829987f",
x"0c998dc998d9",
x"0c998e1998dd",
x"0c998e6998e2",
x"0c9993e9993d",
x"0c9994399941",
x"0c9994899946",
x"0c999a1999a0",
x"0c999a6999a5",
x"0c999ab999aa",
x"0c99a0599a02",
x"0c99a0b99a07",
x"0c99a1099a0c",
x"0c99a1599a11",
x"0c99a6399a60",
x"0c99a6999a65",
x"0c99a6e99a6a",
x"0c99a7499a70",
x"0c99c1799c16",
x"0c99c1a99c18",
x"0c99c7899c74",
x"0c99c7e99c7a",
x"0c99c8399c7f",
x"0c99cdc99cd9",
x"0c99cde99cdd",
x"0c99ce399ce0",
x"0c99ce699ce4",
x"0c99d3e99d3b",
x"0c99d4499d40",
x"0c99d4999d45",
x"0c99da399d9f",
x"0c99da899da4",
x"0c99dad99da9",
x"0c99e0599e03",
x"0c99e0899e06",
x"0c99e0d99e0a",
x"0c99e1299e0f",
x"0c99e1599e14",
x"0c99e6399e62",
x"0c99e6999e67",
x"0c99e6c99e6a",
x"0c99e7199e6d",
x"0c99e7499e72",
x"0c9a0179a015",
x"0c9a01a9a019",
x"0c9a0789a077",
x"0c9a07b9a079",
x"0c9a0809a07c",
x"0c9a0839a081",
x"0c9a0dc9a0d8",
x"0c9a0de9a0dd",
x"0c9a0e39a0e0",
x"0c9a0e69a0e5",
x"0c9a13c9a13b",
x"0c9a1419a13f",
x"0c9a1469a143",
x"0c9a1499a147",
x"0c9a1a09a19e",
x"0c9a1a59a1a1",
x"0c9a1aa9a1a6",
x"0c9a1ad9a1ab",
x"0c9a2059a203",
x"0c9a2089a206",
x"0c9a20d9a20a",
x"0c9a2129a20f",
x"0c9a2159a214",
x"0c9a2639a262",
x"0c9a2699a267",
x"0c9a26c9a26a",
x"0c9a2719a26d",
x"0c9a2749a272",
x"0c9a4179a415",
x"0c9a41a9a419",
x"0c9a4789a476",
x"0c9a47b9a479",
x"0c9a4809a47c",
x"0c9a4839a482",
x"0c9a4d99a4d7",
x"0c9a4de9a4da",
x"0c9a4e39a4e0",
x"0c9a4e69a4e5",
x"0c9a5419a53b",
x"0c9a5469a543",
x"0c9a5499a548",
x"0c9a5a29a59f",
x"0c9a5a59a5a3",
x"0c9a5aa9a5a6",
x"0c9a5ad9a5ac",
x"0c9a6059a603",
x"0c9a6089a606",
x"0c9a60d9a60a",
x"0c9a6129a60f",
x"0c9a6159a614",
x"0c9a6639a662",
x"0c9a6689a666",
x"0c9a66c9a66a",
x"0c9a6719a66d",
x"0c9a6749a672",
x"0c9a8179a816",
x"0c9a81a9a819",
x"0c9a8779a875",
x"0c9a87b9a879",
x"0c9a8809a87c",
x"0c9a8839a881",
x"0c9a8de9a8d7",
x"0c9a8e19a8e0",
x"0c9a8e39a8e2",
x"0c9a8e69a8e4",
x"0c9a93c9a93b",
x"0c9a9419a93d",
x"0c9a9469a943",
x"0c9a9499a948",
x"0c9a9a59a99e",
x"0c9a9aa9a9a6",
x"0c9a9ad9a9ab",
x"0c9aa059aa03",
x"0c9aa0b9aa07",
x"0c9aa109aa0c",
x"0c9aa159aa11",
x"0c9aa649aa61",
x"0c9aa689aa65",
x"0c9aa6c9aa6a",
x"0c9aa719aa6d",
x"0c9aa749aa72",
x"0c9ac1a9ac16",
x"0c9ac789ac74",
x"0c9ac839ac79",
x"0c9acdc9acda",
x"0c9ace19acdd",
x"0c9ace69ace2",
x"0c9ad3c9ad3b",
x"0c9ad419ad3d",
x"0c9ad449ad42",
x"0c9ad469ad45",
x"0c9ad499ad47",
x"0c9ada09ad9e",
x"0c9ada59ada1",
x"0c9adaa9ada6",
x"0c9adad9adab",
x"0c9ae069ae02",
x"0c9ae0b9ae07",
x"0c9ae0f9ae0c",
x"0c9ae159ae11",
x"0c9ae6a9ae60",
x"0c9ae6e9ae6b",
x"0c9ae739ae70",
x"0c9b0189b017",
x"0c9b0799b075",
x"0c9b07d9b07a",
x"0c9b0829b07f",
x"0c9b0e09b0de",
x"0c9b0e59b0e3",
x"0c9b13e9b13b",
x"0c9b1449b140",
x"0c9b1499b145",
x"0c9b1a39b19e",
x"0c9b1a79b1a4",
x"0c9b1ac9b1a9",--fin graph
        x"100000e0146a",                --debut phrase EN217
        x"100001701470",
        x"100000201476",
        x"10000010147c",
        x"100000701482",
        x"100002401488",
        x"10000190148e",
        x"100001b01494",
        x"10000180149a",
        x"100000c014a0",
        x"100000e014a6",
        x"100001c014ac",
        x"100001c014b2",
        x"100000e014b8",
        x"100001e014be",
        x"100001b014c4",
        x"1000024014ca",
        x"1000003014d0",
        x"1000002014d6",
        x"100000b014dc",
        x"1000012014e2",
        x"100001d014e8",
        x"100001c014ee",
        x"1000024014f4",
        x"1000019014fa",
        x"100001801500",
        x"100001e01506",
        x"100001b0150c",
        x"100002401512",
        x"100001501518",
        x"100000e0151e",
        x"100002401524",
        x"100000c0152a",
        x"100000a01530",
        x"100001501536",
        x"100000c0153c",
        x"100001e01542",
        x"100001501548",
        x"10000240154e",
        x"100000d01554",
        x"100000e0155a",
        x"100002401560",
        x"100001701566",
        x"10000180156c",
        x"100001601572",
        x"100000b01578",
        x"100001b0157e",
        x"100000e01584",
        x"100001c0158a",
        x"100002401590",
        x"100001901596",
        x"100001b0159c",
        x"100000e015a2",
        x"1000016015a8",
        x"1000012015ae",
        x"100000e015b4",
        x"100001b015ba",
        x"100001c015c0",                --fin phrase EN217  
        x"100001c64161",
        x"0c1f86b1f86a",                --debut bongo cat
        x"0c1fc6c1fc69",
        x"0c2006d20068",
        x"0c2046e20467",
        x"0c2086f20867",
        x"0c20c7020c66",
        x"0c2107121065",
        x"0c2147221464",
        x"0c2187321863",
        x"0c21c7421c63",
        x"0c2207422062",
        x"0c2247522462",
        x"0c2287722861",
        x"0c22c7a22c60",
        x"0c2307d2305f",
        x"0c234802345c",
        x"0c2388223858",
        x"0c23c8423c55",
        x"0c2408624052",
        x"0c2448824450",
        x"0c2488a2484e",
        x"0c24c8c24c4b",
        x"0c2508d25049",
        x"0c2548f25446",
        x"0c2589025843",
        x"0c25c9225c40",
        x"0c260932603d",
        x"0c264942643b",
        x"0c2689626838",
        x"0c26c9726c36",
        x"0c2709827034",
        x"0c2749a27433",
        x"0c2789b27831",
        x"0c27c9c27c2f",
        x"0c280112800f",
        x"0c2809d2802d",
        x"0c284132840f",
        x"0c2849f2842c",
        x"0c288162880f",
        x"0c288a02882a",
        x"0c28c1828c0f",
        x"0c28ca128c28",
        x"0c2901b2900f",
        x"0c290a229026",
        x"0c2941d2940f",
        x"0c294a329423",
        x"0c2981f2980f",
        x"0c298a429822",
        x"0c29ca529c0f",
        x"0c2a0a62a00f",
        x"0c2a4a82a40f",
        x"0c2a8a82a80f",
        x"0c2ac802ac0f",
        x"0c2aca92ac86",
        x"0c2b07f2b00f",
        x"0c2b0ab2b087",
        x"0c2b47f2b40f",
        x"0c2b4ac2b487",
        x"0c2b87e2b810",
        x"0c2b8ad2b888",
        x"0c2bc7e2bc10",
        x"0c2bcae2bc88",
        x"0c2c07e2c010",
        x"0c2c0af2c088",
        x"0c2c47f2c411",
        x"0c2c4b02c488",
        x"0c2c8762c811",
        x"0c2c87f2c879",
        x"0c2c8b12c888",
        x"0c2cc752cc12",
        x"0c2cc802cc79",
        x"0c2ccb22cc87",
        x"0c2d06b2d012",
        x"0c2d0752d06f",
        x"0c2d0812d079",
        x"0c2d0b22d086",
        x"0c2d46a2d412",
        x"0c2d4b32d479",
        x"0c2d86a2d813",
        x"0c2d8b42d879",
        x"0c2dc6a2dc13",
        x"0c2dcb52dc78",
        x"0c2e0692e013",
        x"0c2e0b52e077",
        x"0c2e4622e413",
        x"0c2e4702e46e",
        x"0c2e4b62e475",
        x"0c2e8612e813",
        x"0c2e8b72e86d",
        x"0c2ec612ec13",
        x"0c2ecb82ec6c",
        x"0c2f0622f014",
        x"0c2f0b92f06b",
        x"0c2f4472f414",
        x"0c2f4b92f44b",
        x"0c2f8462f814",
        x"0c2f8ba2f84d",
        x"0c2fc462fc14",
        x"0c2fcba2fc4e",
        x"0c3004630015",
        x"0c300bb3004e",
        x"0c3044630415",
        x"0c304bb3044e",
        x"0c3084630815",
        x"0c308bb3084f",
        x"0c30c4630c15",
        x"0c30cbb30c4f",
        x"0c3104631014",
        x"0c310923104e",
        x"0c310bb31093",
        x"0c3144731414",
        x"0c314903144e",
        x"0c314bb31496",
        x"0c3184831813",
        x"0c3188b3184b",
        x"0c318bb31899",
        x"0c31c8731c12",
        x"0c31cbb31c9d",
        x"0c3208232011",
        x"0c320bb320a0",
        x"0c3247d32411",
        x"0c324ba324a4",
        x"0c3287832810",
        x"0c328b9328a7",
        x"0c32c7532c10",
        x"0c32cb632ca9",
        x"0c330703300f",
        x"0c3346c3340f",
        x"0c338683380e",
        x"0c33c6433c0e",
        x"0c340453400d",
        x"0c3405f34047",
        x"0c344443440d",
        x"0c3445b34449",
        x"0c348443480c",
        x"0c348573484a",
        x"0c34c4534c0c",
        x"0c34c5334c4b",
        x"0c350463500b",
        x"0c3504e3504b",
        x"0c354473540b",
        x"0c358483580a",
        x"0c35c4935c0a",
        x"0c360493600a",
        x"0c3644a36409",
        x"0c3684b36809",
        x"0c36c4b36c09",
        x"0c3704b37008",
        x"0c3744b37408",
        x"0c3781b37807",
        x"0c3784b37823",
        x"0c37c1a37c07",
        x"0c37c4b37c27",
        x"0c3801a38007",
        x"0c3804b3802a",
        x"0c3841738407",
        x"0c3844b3842d",
        x"0c3881438806",
        x"0c3884b38830",
        x"0c38c1038c06",
        x"0c38c4938c34",
        x"0c3900a39006",
        x"0c3904839037",                --fin bongo cat
        x"0c0046500401",                --debut qr
        x"0c0086500801",
        x"0c00c6500c01",
        x"0c0106501001",
        x"0c0140501401",
        x"0c0142b0141b",
        x"0c014310142e",
        x"0c0143701434",
        x"0c0144a0143b",
        x"0c0146501460",
        x"0c0180501801",
        x"0c0182b0181b",
        x"0c018310182e",
        x"0c0183701834",
        x"0c0184a0183b",
        x"0c0186501860",
        x"0c01c0501c01",
        x"0c01c2b01c1b",
        x"0c01c3101c2e",
        x"0c01c3701c34",
        x"0c01c4a01c3b",
        x"0c01c6501c60",
        x"0c0200502001",
        x"0c0201802009",
        x"0c020210201b",
        x"0c0202702025",
        x"0c0203702034",
        x"0c0203d0203b",
        x"0c0204302041",
        x"0c0204a02047",
        x"0c0205c0204d",
        x"0c0206502060",
        x"0c0240502401",
        x"0c0241802409",
        x"0c024210241b",
        x"0c0242702425",
        x"0c0243702434",
        x"0c0243d0243b",
        x"0c0244302441",
        x"0c0244a02447",
        x"0c0245c0244d",
        x"0c0246502460",
        x"0c0280502801",
        x"0c0281802809",
        x"0c028210281b",
        x"0c0282702825",
        x"0c0283702834",
        x"0c0283d0283b",
        x"0c0284302841",
        x"0c0284a02847",
        x"0c0285c0284d",
        x"0c0286502860",
        x"0c02c0502c01",
        x"0c02c0b02c09",
        x"0c02c1802c15",
        x"0c02c1e02c1b",
        x"0c02c3102c28",
        x"0c02c4a02c3b",
        x"0c02c5002c4d",
        x"0c02c5c02c5a",
        x"0c02c6502c60",
        x"0c0300503001",
        x"0c0300b03009",
        x"0c0301803015",
        x"0c0301e0301b",
        x"0c0303103028",
        x"0c0304a0303b",
        x"0c030500304d",
        x"0c0305c0305a",
        x"0c0306503060",
        x"0c0340503401",
        x"0c0340b03409",
        x"0c0341803415",
        x"0c0341e0341b",
        x"0c0343103428",
        x"0c0344a0343b",
        x"0c034500344d",
        x"0c0345c0345a",
        x"0c0346503460",
        x"0c0380503801",
        x"0c0380b03809",
        x"0c0381803815",
        x"0c038240381b",
        x"0c0383d03837",
        x"0c0384a03847",
        x"0c038500384d",
        x"0c0385c0385a",
        x"0c0386503860",
        x"0c03c0503c01",
        x"0c03c0b03c09",
        x"0c03c1803c15",
        x"0c03c2403c1b",
        x"0c03c3d03c37",
        x"0c03c4a03c47",
        x"0c03c5003c4d",
        x"0c03c5c03c5a",
        x"0c03c6503c60",
        x"0c0400504001",
        x"0c0400b04009",
        x"0c0401804015",
        x"0c040240401b",
        x"0c0403d04037",
        x"0c0404a04047",
        x"0c040500404d",
        x"0c0405c0405a",
        x"0c0406504060",
        x"0c0440504401",
        x"0c0440b04409",
        x"0c0441804415",
        x"0c044240441b",
        x"0c0444a04447",
        x"0c044500444d",
        x"0c0445c0445a",
        x"0c0446504460",
        x"0c0480504801",
        x"0c0480b04809",
        x"0c0481804815",
        x"0c0482e0481b",
        x"0c0483704834",
        x"0c048400483e",
        x"0c0484a04844",
        x"0c048500484d",
        x"0c0485c0485a",
        x"0c0486504860",
        x"0c04c0504c01",
        x"0c04c0b04c09",
        x"0c04c1804c15",
        x"0c04c2e04c1b",
        x"0c04c3704c34",
        x"0c04c4004c3e",
        x"0c04c4a04c44",
        x"0c04c5004c4d",
        x"0c04c5c04c5a",
        x"0c04c6504c60",
        x"0c0500505001",
        x"0c0500c05009",
        x"0c0501805015",
        x"0c0501e0501b",
        x"0c0502705022",
        x"0c050400503e",
        x"0c0504a05047",
        x"0c050500504d",
        x"0c0505c05059",
        x"0c0506505060",
        x"0c0540505401",
        x"0c0541805409",
        x"0c0541e0541b",
        x"0c0542705422",
        x"0c0544005437",
        x"0c0544a05447",
        x"0c0545c0544d",
        x"0c0546505460",
        x"0c0580505801",
        x"0c0581805809",
        x"0c0581e0581b",
        x"0c0582705822",
        x"0c0584005837",
        x"0c0584a05847",
        x"0c0585c0584d",
        x"0c0586505860",
        x"0c05c0505c01",
        x"0c05c1e05c1b",
        x"0c05c2405c22",
        x"0c05c3d05c3b",
        x"0c05c4a05c47",
        x"0c05c6505c60",
        x"0c0600506001",
        x"0c0601e0601b",
        x"0c0602406022",
        x"0c0602b06028",
        x"0c060310602e",
        x"0c0603706034",
        x"0c0603d0603b",
        x"0c0604306041",
        x"0c0604a06047",
        x"0c0606506060",
        x"0c0640506401",
        x"0c0641e0641b",
        x"0c0642406422",
        x"0c0642b06428",
        x"0c064310642e",
        x"0c0643706434",
        x"0c0643d0643b",
        x"0c0644306441",
        x"0c0644a06447",
        x"0c0646506460",
        x"0c0680506801",
        x"0c0681e0681b",
        x"0c0682b06828",
        x"0c068310682e",
        x"0c0683706834",
        x"0c0684a06847",
        x"0c0686506860",
        x"0c06c1e06c01",
        x"0c06c3106c28",
        x"0c06c3a06c34",
        x"0c06c6506c44",
        x"0c0701e07001",
        x"0c0703107028",
        x"0c0703a07034",
        x"0c0706507044",
        x"0c0740807401",
        x"0c0740f0740c",
        x"0c0741507412",
        x"0c0741b07418",
        x"0c0742e07428",
        x"0c0743a07437",
        x"0c074500744d",
        x"0c0746507460",
        x"0c0780807801",
        x"0c0780f0780c",
        x"0c0781507812",
        x"0c0781b07818",
        x"0c0782407822",
        x"0c0782e07828",
        x"0c0784007837",
        x"0c078500784d",
        x"0c0786507860",
        x"0c07c0807c01",
        x"0c07c0f07c0c",
        x"0c07c1507c12",
        x"0c07c1b07c18",
        x"0c07c2407c22",
        x"0c07c2e07c28",
        x"0c07c4007c37",
        x"0c07c5007c4d",
        x"0c07c6507c60",
        x"0c0800808001",
        x"0c0800f0800c",
        x"0c0801b08018",
        x"0c0802e08028",
        x"0c0803d08037",
        x"0c0806508060",
        x"0c0840808401",
        x"0c0840f0840c",
        x"0c0841b08418",
        x"0c0843d08425",
        x"0c0844608441",
        x"0c0844d0844a",
        x"0c0845308450",
        x"0c0845908457",
        x"0c0846508460",
        x"0c0880808801",
        x"0c0880f0880c",
        x"0c0881b08818",
        x"0c0883d08825",
        x"0c0884608841",
        x"0c0884d0884a",
        x"0c0885308850",
        x"0c0885908857",
        x"0c0886508860",
        x"0c08c0808c01",
        x"0c08c0f08c0c",
        x"0c08c1b08c18",
        x"0c08c3d08c25",
        x"0c08c4608c41",
        x"0c08c4d08c4a",
        x"0c08c5308c50",
        x"0c08c5908c57",
        x"0c08c6508c60",
        x"0c0900b09001",
        x"0c0901509012",
        x"0c0902109018",
        x"0c0902709025",
        x"0c0903d0903b",
        x"0c0904609041",
        x"0c090500904d",
        x"0c0905909053",
        x"0c090650905d",
        x"0c0940b09401",
        x"0c0941509412",
        x"0c0942109418",
        x"0c0942709425",
        x"0c0943d0943b",
        x"0c0944609441",
        x"0c094500944d",
        x"0c0945909453",
        x"0c094650945d",
        x"0c0980b09801",
        x"0c0981509812",
        x"0c0982109818",
        x"0c0982709825",
        x"0c0983d0983b",
        x"0c0984609841",
        x"0c098500984d",
        x"0c0985909853",
        x"0c098650985d",
        x"0c09c0509c01",
        x"0c09c0f09c09",
        x"0c09c2109c1f",
        x"0c09c2709c25",
        x"0c09c3409c2b",
        x"0c09c3a09c37",
        x"0c09c4609c3e",
        x"0c09c5009c4a",
        x"0c09c5c09c5a",
        x"0c09c6509c60",
        x"0c0a0050a001",
        x"0c0a00f0a009",
        x"0c0a0210a01f",
        x"0c0a0270a025",
        x"0c0a0340a02b",
        x"0c0a03a0a037",
        x"0c0a0460a03e",
        x"0c0a0500a04a",
        x"0c0a05c0a05a",
        x"0c0a0650a060",
        x"0c0a4050a401",
        x"0c0a40f0a409",
        x"0c0a4210a41f",
        x"0c0a4270a425",
        x"0c0a4340a42b",
        x"0c0a43a0a437",
        x"0c0a4460a43e",
        x"0c0a4500a44a",
        x"0c0a45c0a45a",
        x"0c0a4650a460",
        x"0c0a8120a801",
        x"0c0a8240a822",
        x"0c0a82e0a82b",
        x"0c0a83d0a831",
        x"0c0a8560a84d",
        x"0c0a8650a85d",
        x"0c0ac120ac01",
        x"0c0ac240ac22",
        x"0c0ac2e0ac2b",
        x"0c0ac3d0ac31",
        x"0c0ac560ac4d",
        x"0c0ac650ac5d",
        x"0c0b0120b001",
        x"0c0b0240b022",
        x"0c0b02e0b02b",
        x"0c0b03d0b031",
        x"0c0b0560b04d",
        x"0c0b0650b05d",
        x"0c0b4080b401",
        x"0c0b40f0b40c",
        x"0c0b41b0b412",
        x"0c0b4240b422",
        x"0c0b42b0b428",
        x"0c0b4370b42e",
        x"0c0b4430b43e",
        x"0c0b44d0b447",
        x"0c0b4590b453",
        x"0c0b4650b460",
        x"0c0b8080b801",
        x"0c0b80f0b80c",
        x"0c0b81b0b812",
        x"0c0b8240b822",
        x"0c0b82b0b828",
        x"0c0b8370b82e",
        x"0c0b8430b83e",
        x"0c0b84d0b847",
        x"0c0b8590b853",
        x"0c0b8650b860",
        x"0c0bc080bc01",
        x"0c0bc0f0bc0c",
        x"0c0bc1b0bc12",
        x"0c0bc240bc22",
        x"0c0bc2b0bc28",
        x"0c0bc370bc2e",
        x"0c0bc430bc3e",
        x"0c0bc4d0bc47",
        x"0c0bc590bc53",
        x"0c0bc650bc60",
        x"0c0c0050c001",
        x"0c0c0210c012",
        x"0c0c0270c025",
        x"0c0c0310c02b",
        x"0c0c03d0c03b",
        x"0c0c04a0c047",
        x"0c0c0650c060",
        x"0c0c4050c401",
        x"0c0c4210c412",
        x"0c0c4270c425",
        x"0c0c4310c42b",
        x"0c0c43d0c43b",
        x"0c0c44a0c447",
        x"0c0c4650c460",
        x"0c0c8050c801",
        x"0c0c8210c812",
        x"0c0c8270c825",
        x"0c0c8310c82b",
        x"0c0c83d0c83b",
        x"0c0c84a0c847",
        x"0c0c8650c860",
        x"0c0cc050cc01",
        x"0c0cc1e0cc1b",
        x"0c0cc650cc60",
        x"0c0d0050d001",
        x"0c0d0120d00c",
        x"0c0d01e0d01b",
        x"0c0d02b0d028",
        x"0c0d03a0d031",
        x"0c0d0400d03e",
        x"0c0d04d0d04a",
        x"0c0d0590d050",
        x"0c0d0650d05d",
        x"0c0d4050d401",
        x"0c0d4120d40c",
        x"0c0d41e0d41b",
        x"0c0d42b0d428",
        x"0c0d43a0d431",
        x"0c0d4400d43e",
        x"0c0d44d0d44a",
        x"0c0d4590d450",
        x"0c0d4650d45d",
        x"0c0d8050d801",
        x"0c0d8120d80c",
        x"0c0d81e0d81b",
        x"0c0d82b0d828",
        x"0c0d8370d834",
        x"0c0d8590d853",
        x"0c0d8650d85d",
        x"0c0dc150dc01",
        x"0c0dc1e0dc18",
        x"0c0dc2b0dc22",
        x"0c0dc370dc34",
        x"0c0dc3d0dc3b",
        x"0c0dc460dc41",
        x"0c0dc650dc53",
        x"0c0e0150e001",
        x"0c0e01e0e018",
        x"0c0e02b0e022",
        x"0c0e0370e034",
        x"0c0e03d0e03b",
        x"0c0e0460e041",
        x"0c0e0650e053",
        x"0c0e4080e401",
        x"0c0e40f0e40c",
        x"0c0e41e0e418",
        x"0c0e42b0e425",
        x"0c0e4370e434",
        x"0c0e4460e441",
        x"0c0e4560e453",
        x"0c0e4650e460",
        x"0c0e8080e801",
        x"0c0e80f0e80c",
        x"0c0e81e0e818",
        x"0c0e82b0e825",
        x"0c0e8370e831",
        x"0c0e8560e83e",
        x"0c0e8650e860",
        x"0c0ec080ec01",
        x"0c0ec0f0ec0c",
        x"0c0ec1e0ec18",
        x"0c0ec2b0ec25",
        x"0c0ec370ec31",
        x"0c0ec560ec3e",
        x"0c0ec650ec60",
        x"0c0f0080f001",
        x"0c0f01e0f018",
        x"0c0f0270f025",
        x"0c0f0460f044",
        x"0c0f0500f04d",
        x"0c0f0650f060",
        x"0c0f4080f401",
        x"0c0f4210f412",
        x"0c0f4270f425",
        x"0c0f42e0f42b",
        x"0c0f43d0f437",
        x"0c0f4460f444",
        x"0c0f4500f44d",
        x"0c0f45c0f45a",
        x"0c0f4650f460",
        x"0c0f8080f801",
        x"0c0f8210f812",
        x"0c0f8270f825",
        x"0c0f82e0f82b",
        x"0c0f83d0f837",
        x"0c0f8460f844",
        x"0c0f8500f84d",
        x"0c0f85c0f85a",
        x"0c0f8650f860",
        x"0c0fc050fc01",
        x"0c0fc3a0fc37",
        x"0c0fc460fc44",
        x"0c0fc500fc4d",
        x"0c0fc5c0fc5a",
        x"0c0fc650fc60",
        x"0c1000510001",
        x"0c1001210009",
        x"0c1003410031",
        x"0c1003a10037",
        x"0c1005310041",
        x"0c1005c1005a",
        x"0c1006510060",
        x"0c1040510401",
        x"0c1041210409",
        x"0c1043410431",
        x"0c1043a10437",
        x"0c1045310441",
        x"0c1045c1045a",
        x"0c1046510460",
        x"0c1080510801",
        x"0c1083a10837",
        x"0c1084310841",
        x"0c1084a10847",
        x"0c108531084d",
        x"0c1085c1085a",
        x"0c1086510860",
        x"0c10c0810c01",
        x"0c10c2710c22",
        x"0c10c4310c34",
        x"0c10c4a10c47",
        x"0c10c5310c4d",
        x"0c10c5c10c57",
        x"0c10c6510c60",
        x"0c1100811001",
        x"0c1102711022",
        x"0c1104311034",
        x"0c1104a11047",
        x"0c110531104d",
        x"0c1105c11057",
        x"0c1106511060",
        x"0c1140811401",
        x"0c1142711422",
        x"0c1144311434",
        x"0c1144a11447",
        x"0c114531144d",
        x"0c1145c11457",
        x"0c1146511460",
        x"0c1180811801",
        x"0c118121180c",
        x"0c1181e11815",
        x"0c1182b11828",
        x"0c1183d1182e",
        x"0c1186511847",
        x"0c11c0811c01",
        x"0c11c1211c0c",
        x"0c11c1e11c15",
        x"0c11c2b11c28",
        x"0c11c3d11c2e",
        x"0c11c6511c47",
        x"0c1200812001",
        x"0c120121200c",
        x"0c1201e12015",
        x"0c1202b12028",
        x"0c1203d1202e",
        x"0c1206512047",
        x"0c1240b12401",
        x"0c1241812415",
        x"0c1241e1241b",
        x"0c1242712425",
        x"0c124311242b",
        x"0c1244312434",
        x"0c1244a12447",
        x"0c1246512460",
        x"0c1280b12801",
        x"0c1281812815",
        x"0c1281e1281b",
        x"0c1282712825",
        x"0c128311282b",
        x"0c1284312834",
        x"0c1284a12847",
        x"0c1286512860",
        x"0c12c0b12c01",
        x"0c12c1812c15",
        x"0c12c1e12c1b",
        x"0c12c2712c25",
        x"0c12c3112c2b",
        x"0c12c4312c34",
        x"0c12c4a12c47",
        x"0c12c6512c60",
        x"0c1300513001",
        x"0c130121300f",
        x"0c1301e13015",
        x"0c1302413022",
        x"0c1303113028",
        x"0c1303a13037",
        x"0c1304a13044",
        x"0c1305c1304d",
        x"0c1306513060",
        x"0c1340513401",
        x"0c134121340f",
        x"0c1341e13415",
        x"0c1342413422",
        x"0c1343113428",
        x"0c1343a13437",
        x"0c1344a13444",
        x"0c1345c1344d",
        x"0c1346513460",
        x"0c1380513801",
        x"0c138121380f",
        x"0c1381e13815",
        x"0c1382413822",
        x"0c1383113828",
        x"0c1383a13837",
        x"0c1384a13844",
        x"0c1385c1384d",
        x"0c1386513860",
        x"0c13c0513c01",
        x"0c13c1213c0f",
        x"0c13c2413c22",
        x"0c13c2b13c28",
        x"0c13c4313c37",
        x"0c13c4a13c47",
        x"0c13c5013c4d",
        x"0c13c5c13c5a",
        x"0c13c6513c60",
        x"0c1400514001",
        x"0c140121400f",
        x"0c1402414022",
        x"0c1402b14028",
        x"0c1404314037",
        x"0c1404a14047",
        x"0c140501404d",
        x"0c1405c1405a",
        x"0c1406514060",
        x"0c1440514401",
        x"0c144121440f",
        x"0c1442414422",
        x"0c1442b14428",
        x"0c1444314437",
        x"0c1444a14447",
        x"0c144501444d",
        x"0c1445c1445a",
        x"0c1446514460",
        x"0c1481514801",
        x"0c1481b14818",
        x"0c1482b14822",
        x"0c1483a14834",
        x"0c148431483e",
        x"0c1484a14847",
        x"0c148501484d",
        x"0c1485c1485a",
        x"0c1486514860",
        x"0c14c1514c01",
        x"0c14c1b14c18",
        x"0c14c2b14c22",
        x"0c14c3a14c34",
        x"0c14c4314c3e",
        x"0c14c4a14c47",
        x"0c14c5014c4d",
        x"0c14c5c14c5a",
        x"0c14c6514c60",
        x"0c1501515001",
        x"0c1501b15018",
        x"0c1502b15022",
        x"0c1503a15034",
        x"0c150431503e",
        x"0c1504a15047",
        x"0c150501504d",
        x"0c1505c1505a",
        x"0c1506515060",
        x"0c1540815401",
        x"0c154151540f",
        x"0c1542715425",
        x"0c1544a15447",
        x"0c154501544d",
        x"0c1545c1545a",
        x"0c1546515460",
        x"0c1580815801",
        x"0c158151580f",
        x"0c158211581f",
        x"0c1582715825",
        x"0c1582e1582b",
        x"0c1584a15847",
        x"0c158501584d",
        x"0c1585c1585a",
        x"0c1586515860",
        x"0c15c0815c01",
        x"0c15c1515c0f",
        x"0c15c2115c1f",
        x"0c15c2715c25",
        x"0c15c2e15c2b",
        x"0c15c4a15c47",
        x"0c15c5015c4d",
        x"0c15c5c15c5a",
        x"0c15c6515c60",
        x"0c1600516001",
        x"0c1601516012",
        x"0c1602716025",
        x"0c1604a16047",
        x"0c160501604d",
        x"0c1605c16059",
        x"0c1606516060",
        x"0c1640516401",
        x"0c1640b16409",
        x"0c1641b16412",
        x"0c1642b16422",
        x"0c164311642e",
        x"0c1643a16434",
        x"0c1644316441",
        x"0c1644a16447",
        x"0c1645c1644d",
        x"0c1646516460",
        x"0c1680516801",
        x"0c1680b16809",
        x"0c1681b16812",
        x"0c1682b16822",
        x"0c168311682e",
        x"0c1683a16834",
        x"0c1684316841",
        x"0c1684a16847",
        x"0c1685c1684d",
        x"0c1686516860",
        x"0c16c0516c01",
        x"0c16c0b16c09",
        x"0c16c1816c15",
        x"0c16c2716c25",
        x"0c16c3a16c37",
        x"0c16c4a16c47",
        x"0c16c6516c60",
        x"0c1700b17001",
        x"0c1701817015",
        x"0c1702717025",
        x"0c1702e1702b",
        x"0c1703417031",
        x"0c1704017037",
        x"0c1704a17047",
        x"0c1706517060",
        x"0c1740b17401",
        x"0c1741817415",
        x"0c1742717425",
        x"0c1742e1742b",
        x"0c1743417431",
        x"0c1744017437",
        x"0c1744a17447",
        x"0c1746517460",
        x"0c1780b17801",
        x"0c1781817815",
        x"0c1782717825",
        x"0c1782e1782b",
        x"0c1783417831",
        x"0c1784017837",
        x"0c1784a17847",
        x"0c1786517860",
        x"0c17c6517c01",
        x"0c1806518001",                --fin qr

        OTHERS => x"000000000000");
BEGIN

    PROCESS(clk)
    BEGIN
        IF falling_edge(clk) THEN
            IF ce = '1' THEN
                data_out_read_only <= memory_data(to_integer(unsigned(address_read_only)));
                IF rw = '1' THEN        -- write
                    memory_data(to_integer(unsigned(address))) <= input;
                ELSE                    --read
                    data_out <= memory_data(to_integer(unsigned(address)));
                END IF;
            END IF;
        END IF;
    END PROCESS;

END Behavioral;
