----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06.02.2023 09:11:07
-- Design Name: 
-- Module Name: glyph_memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY glyph_memory IS
    PORT (
        clk : IN STD_LOGIC;
        ce : IN STD_LOGIC;
        number : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
        data_out : OUT STD_LOGIC_VECTOR(39 DOWNTO 0));
END glyph_memory;

ARCHITECTURE Behavioral OF glyph_memory IS
    TYPE memory_array IS ARRAY (INTEGER RANGE 0 TO 63) OF STD_LOGIC_VECTOR (39 DOWNTO 0);
    SIGNAL memory_data : memory_array := (
        "0111010001100011000110001100011000101110", --0
        "0010001100101000010000100001000010011111", --1
        "0111010001000010000100010001000100011111", --2
        "0111010001000010000100111000011000101110", --3
        "0001000100010001010011111001000010000100", --4
        "1111110000100001111000001000010000101110", --5
        "0111010000100001111010001100011000101110", --6
        "1111100001000100010001000100001000010000", --7
        "0111010001100010111010001100011000101110", --8
        "0111010001100011000101111000010000101110", --9
        "0111010001100011000111111100011000110001", --A
        "1111010001100011111110001100011000111110", --B
        "0111110000100001000010000100001000001111", --C
        "1111010001100011000110001100011000111110", --D
        "1111110000100001000011100100001000011111", --E
        "1111110000100001110010000100001000010000", --F
        "0111010001100001000010111100011000101110", --G
        "1000110001100011000111111100011000110001", --H
        "0000000100000000010000100001000010000100", --I
        "0111000100001000010000100101001010001000", --J
        "1000010001100101010011000101001001010001", --K
        "1000010000100001000010000100001000011111", --L
        "1000111011101011000110001100011000110001", --M
        "1000110001110011010110101100111000110001", --N
        "0111010001100011000110001100011000101110", --0
        "0111010001100011000111110100001000010000", --P
        "0111010001100011000110001101011001001101", --Q
        "0111010001100011000111110101001001010001", --R
        "0111110000100001000001110000010000111110", --S
        "1111100100001000010000100001000010000100", --T
        "1000110001100011000110001100011000101110", --U
        "1000110001100011000110001100010101000100", --V
        "1000110001100011000110001100011010101010", --W
        "1000110001010100010001010100011000110001", --X
        "1000110001010100010000100001000010000100", --Y
        "1111100001000010001000100010001000011111", --Z  
        "0000000000000000000000000000000000000000", --VIDE
        OTHERS => "1111111111111111111111111111111111111111");
BEGIN

    PROCESS (clk)
    BEGIN
        IF falling_edge(clk) THEN
            IF ce = '1' THEN
                data_out <= memory_data(to_integer(unsigned(number)));
            END IF;
        END IF;
    END PROCESS;

END Behavioral;